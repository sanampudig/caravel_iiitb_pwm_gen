magic
tech sky130B
magscale 1 2
timestamp 1662984762
<< obsli1 >>
rect 1104 2159 28888 27761
<< obsm1 >>
rect 14 2128 28888 27792
<< metal2 >>
rect 18050 29200 18106 30000
rect 18 0 74 800
rect 23202 0 23258 800
<< obsm2 >>
rect 20 29144 17994 29200
rect 18162 29144 28226 29200
rect 20 856 28226 29144
rect 130 800 23146 856
rect 23314 800 28226 856
<< metal3 >>
rect 0 24488 800 24608
rect 29200 17008 30000 17128
<< obsm3 >>
rect 800 24688 29200 27777
rect 880 24408 29200 24688
rect 800 17208 29200 24408
rect 800 16928 29120 17208
rect 800 2143 29200 16928
<< metal4 >>
rect 4418 2128 4738 27792
rect 7892 2128 8212 27792
rect 11366 2128 11686 27792
rect 14840 2128 15160 27792
rect 18314 2128 18634 27792
rect 21788 2128 22108 27792
rect 25262 2128 25582 27792
<< labels >>
rlabel metal3 s 0 24488 800 24608 6 PWM_OUT
port 1 nsew signal output
rlabel metal2 s 18 0 74 800 6 clk
port 2 nsew signal input
rlabel metal3 s 29200 17008 30000 17128 6 decrease_duty
port 3 nsew signal input
rlabel metal2 s 18050 29200 18106 30000 6 increase_duty
port 4 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 reset
port 5 nsew signal input
rlabel metal4 s 4418 2128 4738 27792 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 11366 2128 11686 27792 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 18314 2128 18634 27792 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 25262 2128 25582 27792 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 7892 2128 8212 27792 6 vssd1
port 7 nsew ground bidirectional
rlabel metal4 s 14840 2128 15160 27792 6 vssd1
port 7 nsew ground bidirectional
rlabel metal4 s 21788 2128 22108 27792 6 vssd1
port 7 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 893376
string GDS_FILE /home/parallels/Desktop/caravel_iiitb_pwm_gen/openlane/iiitb_pwm_gen/runs/22_09_12_17_41/results/signoff/iiitb_pwm_gen.magic.gds
string GDS_START 257440
<< end >>

