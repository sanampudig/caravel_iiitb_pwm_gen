magic
tech sky130B
magscale 1 2
timestamp 1662984761
<< viali >>
rect 17693 27557 17727 27591
rect 18337 27421 18371 27455
rect 18153 27285 18187 27319
rect 1685 24769 1719 24803
rect 1501 24565 1535 24599
rect 3525 20417 3559 20451
rect 3433 20213 3467 20247
rect 3985 20213 4019 20247
rect 2789 19805 2823 19839
rect 3801 19805 3835 19839
rect 2881 19669 2915 19703
rect 4997 17221 5031 17255
rect 4813 17153 4847 17187
rect 5089 17153 5123 17187
rect 7849 17153 7883 17187
rect 8953 17153 8987 17187
rect 27537 17153 27571 17187
rect 28181 17153 28215 17187
rect 7941 17085 7975 17119
rect 9045 17085 9079 17119
rect 7481 17017 7515 17051
rect 8585 17017 8619 17051
rect 4629 16949 4663 16983
rect 27997 16949 28031 16983
rect 9137 16745 9171 16779
rect 5089 16609 5123 16643
rect 7757 16609 7791 16643
rect 8217 16609 8251 16643
rect 10517 16609 10551 16643
rect 11345 16609 11379 16643
rect 4813 16541 4847 16575
rect 4997 16541 5031 16575
rect 5181 16541 5215 16575
rect 5365 16541 5399 16575
rect 7113 16541 7147 16575
rect 8125 16541 8159 16575
rect 9321 16541 9355 16575
rect 9413 16541 9447 16575
rect 9597 16541 9631 16575
rect 9689 16541 9723 16575
rect 10149 16541 10183 16575
rect 10333 16541 10367 16575
rect 11529 16541 11563 16575
rect 11805 16541 11839 16575
rect 5549 16405 5583 16439
rect 7021 16405 7055 16439
rect 11713 16405 11747 16439
rect 4721 16201 4755 16235
rect 7849 16201 7883 16235
rect 9321 16201 9355 16235
rect 6377 16133 6411 16167
rect 4905 16065 4939 16099
rect 4997 16065 5031 16099
rect 5273 16065 5307 16099
rect 6561 16065 6595 16099
rect 6653 16065 6687 16099
rect 8953 16065 8987 16099
rect 11713 16065 11747 16099
rect 3617 15997 3651 16031
rect 3893 15997 3927 16031
rect 5181 15997 5215 16031
rect 7941 15997 7975 16031
rect 8125 15997 8159 16031
rect 9045 15997 9079 16031
rect 6377 15929 6411 15963
rect 7481 15861 7515 15895
rect 11805 15861 11839 15895
rect 12173 15861 12207 15895
rect 7389 15657 7423 15691
rect 9229 15589 9263 15623
rect 5365 15521 5399 15555
rect 6561 15521 6595 15555
rect 8953 15521 8987 15555
rect 13369 15521 13403 15555
rect 5733 15453 5767 15487
rect 5825 15453 5859 15487
rect 6653 15453 6687 15487
rect 7481 15453 7515 15487
rect 9137 15453 9171 15487
rect 9321 15453 9355 15487
rect 9413 15453 9447 15487
rect 11345 15453 11379 15487
rect 12081 15453 12115 15487
rect 6009 15385 6043 15419
rect 5457 15317 5491 15351
rect 5641 15317 5675 15351
rect 11897 15317 11931 15351
rect 12817 15317 12851 15351
rect 13185 15317 13219 15351
rect 13277 15317 13311 15351
rect 4905 15113 4939 15147
rect 6469 15113 6503 15147
rect 12633 15113 12667 15147
rect 4537 15045 4571 15079
rect 2145 14977 2179 15011
rect 2329 14977 2363 15011
rect 4445 14977 4479 15011
rect 4721 14977 4755 15011
rect 6561 14977 6595 15011
rect 12265 14977 12299 15011
rect 12173 14909 12207 14943
rect 2145 14773 2179 14807
rect 7757 14773 7791 14807
rect 7389 14569 7423 14603
rect 11805 14569 11839 14603
rect 2513 14501 2547 14535
rect 4077 14501 4111 14535
rect 11529 14433 11563 14467
rect 2329 14365 2363 14399
rect 2605 14365 2639 14399
rect 3249 14365 3283 14399
rect 3801 14365 3835 14399
rect 4077 14365 4111 14399
rect 5181 14365 5215 14399
rect 6653 14365 6687 14399
rect 7297 14365 7331 14399
rect 7573 14365 7607 14399
rect 8401 14365 8435 14399
rect 10701 14365 10735 14399
rect 10793 14365 10827 14399
rect 11345 14365 11379 14399
rect 11437 14365 11471 14399
rect 11621 14365 11655 14399
rect 12449 14365 12483 14399
rect 8309 14297 8343 14331
rect 9873 14297 9907 14331
rect 12357 14297 12391 14331
rect 2145 14229 2179 14263
rect 3065 14229 3099 14263
rect 3893 14229 3927 14263
rect 5089 14229 5123 14263
rect 6469 14229 6503 14263
rect 7757 14229 7791 14263
rect 9781 14229 9815 14263
rect 2145 14025 2179 14059
rect 7205 14025 7239 14059
rect 8769 14025 8803 14059
rect 10333 14025 10367 14059
rect 13001 14025 13035 14059
rect 9873 13957 9907 13991
rect 13461 13957 13495 13991
rect 2789 13889 2823 13923
rect 2881 13889 2915 13923
rect 3065 13889 3099 13923
rect 3893 13889 3927 13923
rect 5457 13889 5491 13923
rect 8033 13889 8067 13923
rect 8125 13889 8159 13923
rect 8953 13889 8987 13923
rect 9229 13889 9263 13923
rect 10149 13889 10183 13923
rect 13185 13889 13219 13923
rect 14013 13889 14047 13923
rect 14105 13889 14139 13923
rect 1685 13821 1719 13855
rect 2605 13821 2639 13855
rect 3617 13821 3651 13855
rect 5365 13821 5399 13855
rect 7021 13821 7055 13855
rect 7113 13821 7147 13855
rect 9965 13821 9999 13855
rect 12265 13821 12299 13855
rect 12541 13821 12575 13855
rect 13369 13821 13403 13855
rect 1961 13753 1995 13787
rect 2973 13753 3007 13787
rect 5825 13753 5859 13787
rect 9045 13753 9079 13787
rect 9137 13753 9171 13787
rect 7573 13685 7607 13719
rect 10149 13685 10183 13719
rect 13277 13685 13311 13719
rect 2329 13481 2363 13515
rect 10517 13481 10551 13515
rect 10701 13481 10735 13515
rect 14105 13481 14139 13515
rect 14473 13481 14507 13515
rect 15025 13413 15059 13447
rect 2697 13345 2731 13379
rect 2789 13345 2823 13379
rect 6653 13345 6687 13379
rect 6837 13345 6871 13379
rect 10793 13345 10827 13379
rect 12541 13345 12575 13379
rect 1685 13277 1719 13311
rect 1869 13277 1903 13311
rect 2513 13277 2547 13311
rect 2605 13277 2639 13311
rect 4445 13277 4479 13311
rect 5089 13277 5123 13311
rect 5733 13277 5767 13311
rect 7941 13277 7975 13311
rect 9045 13277 9079 13311
rect 9689 13277 9723 13311
rect 10057 13277 10091 13311
rect 10885 13277 10919 13311
rect 11529 13277 11563 13311
rect 14381 13277 14415 13311
rect 14473 13277 14507 13311
rect 15209 13277 15243 13311
rect 4261 13209 4295 13243
rect 9873 13209 9907 13243
rect 12449 13209 12483 13243
rect 1777 13141 1811 13175
rect 4997 13141 5031 13175
rect 5641 13141 5675 13175
rect 6193 13141 6227 13175
rect 6561 13141 6595 13175
rect 7849 13141 7883 13175
rect 9137 13141 9171 13175
rect 11345 13141 11379 13175
rect 11989 13141 12023 13175
rect 12357 13141 12391 13175
rect 2237 12937 2271 12971
rect 3709 12937 3743 12971
rect 14749 12937 14783 12971
rect 2145 12801 2179 12835
rect 2421 12801 2455 12835
rect 4353 12801 4387 12835
rect 4997 12801 5031 12835
rect 5457 12801 5491 12835
rect 7021 12801 7055 12835
rect 7481 12801 7515 12835
rect 9413 12801 9447 12835
rect 11989 12801 12023 12835
rect 14105 12801 14139 12835
rect 14565 12801 14599 12835
rect 4905 12733 4939 12767
rect 13829 12733 13863 12767
rect 2421 12665 2455 12699
rect 5549 12665 5583 12699
rect 14013 12665 14047 12699
rect 4261 12597 4295 12631
rect 6929 12597 6963 12631
rect 7665 12597 7699 12631
rect 9505 12597 9539 12631
rect 11805 12597 11839 12631
rect 13921 12597 13955 12631
rect 15393 12393 15427 12427
rect 14197 12257 14231 12291
rect 5181 12189 5215 12223
rect 14381 12189 14415 12223
rect 14473 12189 14507 12223
rect 4997 12053 5031 12087
rect 14841 12053 14875 12087
rect 9597 11849 9631 11883
rect 7849 11645 7883 11679
rect 8125 11645 8159 11679
rect 4629 11509 4663 11543
rect 10701 11509 10735 11543
rect 11713 11509 11747 11543
rect 3249 11305 3283 11339
rect 5733 11305 5767 11339
rect 12265 11305 12299 11339
rect 14841 11305 14875 11339
rect 1777 11169 1811 11203
rect 4261 11169 4295 11203
rect 10793 11169 10827 11203
rect 1501 11101 1535 11135
rect 3985 11101 4019 11135
rect 10517 11101 10551 11135
rect 14749 11101 14783 11135
rect 9045 10761 9079 10795
rect 13277 10761 13311 10795
rect 2145 10693 2179 10727
rect 4353 10693 4387 10727
rect 10517 10693 10551 10727
rect 1869 10625 1903 10659
rect 6745 10625 6779 10659
rect 15025 10625 15059 10659
rect 4077 10557 4111 10591
rect 6377 10557 6411 10591
rect 8217 10557 8251 10591
rect 10793 10557 10827 10591
rect 11529 10557 11563 10591
rect 11805 10557 11839 10591
rect 14841 10489 14875 10523
rect 3617 10421 3651 10455
rect 5825 10421 5859 10455
rect 3249 10217 3283 10251
rect 7987 10149 8021 10183
rect 1777 10081 1811 10115
rect 6193 10081 6227 10115
rect 6561 10081 6595 10115
rect 10609 10081 10643 10115
rect 14565 10081 14599 10115
rect 1501 10013 1535 10047
rect 10333 10013 10367 10047
rect 14657 10013 14691 10047
rect 12081 9877 12115 9911
rect 2053 9605 2087 9639
rect 11805 9605 11839 9639
rect 8401 9537 8435 9571
rect 11529 9537 11563 9571
rect 14013 9537 14047 9571
rect 14105 9537 14139 9571
rect 15301 9537 15335 9571
rect 19073 9537 19107 9571
rect 19533 9537 19567 9571
rect 1777 9469 1811 9503
rect 3525 9469 3559 9503
rect 6653 9469 6687 9503
rect 8125 9469 8159 9503
rect 13277 9469 13311 9503
rect 15025 9469 15059 9503
rect 14013 9333 14047 9367
rect 14381 9333 14415 9367
rect 16681 9333 16715 9367
rect 18981 9333 19015 9367
rect 19625 9333 19659 9367
rect 7757 9129 7791 9163
rect 14381 9129 14415 9163
rect 6009 8993 6043 9027
rect 10057 8925 10091 8959
rect 14473 8925 14507 8959
rect 6285 8857 6319 8891
rect 9505 8517 9539 8551
rect 3249 8449 3283 8483
rect 9229 8449 9263 8483
rect 14105 8449 14139 8483
rect 3525 8381 3559 8415
rect 14013 8381 14047 8415
rect 4997 8313 5031 8347
rect 7113 8313 7147 8347
rect 10977 8313 11011 8347
rect 11529 8245 11563 8279
rect 3801 8041 3835 8075
rect 9781 8041 9815 8075
rect 13461 8041 13495 8075
rect 14105 8041 14139 8075
rect 14565 8041 14599 8075
rect 15209 8041 15243 8075
rect 15577 8041 15611 8075
rect 1501 7905 1535 7939
rect 8401 7905 8435 7939
rect 10609 7905 10643 7939
rect 10885 7905 10919 7939
rect 14197 7905 14231 7939
rect 13553 7837 13587 7871
rect 14381 7837 14415 7871
rect 15209 7837 15243 7871
rect 15393 7837 15427 7871
rect 1777 7769 1811 7803
rect 6653 7769 6687 7803
rect 14105 7769 14139 7803
rect 16497 7769 16531 7803
rect 16681 7769 16715 7803
rect 3249 7701 3283 7735
rect 6193 7701 6227 7735
rect 12357 7701 12391 7735
rect 17325 7701 17359 7735
rect 3065 7497 3099 7531
rect 10977 7497 11011 7531
rect 14105 7497 14139 7531
rect 6745 7429 6779 7463
rect 1961 7361 1995 7395
rect 4353 7361 4387 7395
rect 9229 7361 9263 7395
rect 13553 7361 13587 7395
rect 14197 7361 14231 7395
rect 14841 7361 14875 7395
rect 9505 7293 9539 7327
rect 13461 7225 13495 7259
rect 4997 7157 5031 7191
rect 5825 7157 5859 7191
rect 8033 7157 8067 7191
rect 14749 7157 14783 7191
rect 4432 6953 4466 6987
rect 6634 6953 6668 6987
rect 14105 6953 14139 6987
rect 4169 6817 4203 6851
rect 14197 6817 14231 6851
rect 2329 6749 2363 6783
rect 3157 6749 3191 6783
rect 6377 6749 6411 6783
rect 10885 6749 10919 6783
rect 14381 6749 14415 6783
rect 16497 6749 16531 6783
rect 1869 6681 1903 6715
rect 11161 6681 11195 6715
rect 14105 6681 14139 6715
rect 3065 6613 3099 6647
rect 5917 6613 5951 6647
rect 8125 6613 8159 6647
rect 12633 6613 12667 6647
rect 14565 6613 14599 6647
rect 16589 6613 16623 6647
rect 4721 6409 4755 6443
rect 8125 6409 8159 6443
rect 13277 6409 13311 6443
rect 14197 6409 14231 6443
rect 14841 6409 14875 6443
rect 2329 6341 2363 6375
rect 5365 6341 5399 6375
rect 6653 6341 6687 6375
rect 12817 6341 12851 6375
rect 4813 6273 4847 6307
rect 11529 6273 11563 6307
rect 13093 6273 13127 6307
rect 13737 6273 13771 6307
rect 14013 6273 14047 6307
rect 14657 6273 14691 6307
rect 2053 6205 2087 6239
rect 6377 6205 6411 6239
rect 8585 6205 8619 6239
rect 8861 6205 8895 6239
rect 10333 6205 10367 6239
rect 12909 6205 12943 6239
rect 13829 6205 13863 6239
rect 3801 6069 3835 6103
rect 12817 6069 12851 6103
rect 14013 6069 14047 6103
rect 6377 5865 6411 5899
rect 6837 5865 6871 5899
rect 8953 5865 8987 5899
rect 11437 5865 11471 5899
rect 13461 5797 13495 5831
rect 6561 5729 6595 5763
rect 9689 5729 9723 5763
rect 16037 5729 16071 5763
rect 6377 5661 6411 5695
rect 6653 5661 6687 5695
rect 13553 5661 13587 5695
rect 14381 5661 14415 5695
rect 15117 5661 15151 5695
rect 15945 5661 15979 5695
rect 9965 5593 9999 5627
rect 14197 5525 14231 5559
rect 14933 5525 14967 5559
rect 9137 5321 9171 5355
rect 7849 5253 7883 5287
rect 4997 5185 5031 5219
rect 5273 5185 5307 5219
rect 10057 5185 10091 5219
rect 13829 5185 13863 5219
rect 2789 5117 2823 5151
rect 3065 5117 3099 5151
rect 4537 5117 4571 5151
rect 5089 5117 5123 5151
rect 5457 5049 5491 5083
rect 2145 4981 2179 5015
rect 4997 4981 5031 5015
rect 6745 4981 6779 5015
rect 11713 4981 11747 5015
rect 13737 4981 13771 5015
rect 3801 4777 3835 4811
rect 8125 4777 8159 4811
rect 13461 4777 13495 4811
rect 16957 4777 16991 4811
rect 19901 4777 19935 4811
rect 3249 4709 3283 4743
rect 12081 4709 12115 4743
rect 1501 4641 1535 4675
rect 6377 4641 6411 4675
rect 6653 4641 6687 4675
rect 10333 4641 10367 4675
rect 14197 4641 14231 4675
rect 4721 4573 4755 4607
rect 13553 4573 13587 4607
rect 14289 4573 14323 4607
rect 14933 4573 14967 4607
rect 16497 4573 16531 4607
rect 19809 4573 19843 4607
rect 1777 4505 1811 4539
rect 10609 4505 10643 4539
rect 14841 4505 14875 4539
rect 4629 4437 4663 4471
rect 16405 4437 16439 4471
rect 11805 4165 11839 4199
rect 6377 4097 6411 4131
rect 11529 4097 11563 4131
rect 2053 4029 2087 4063
rect 2329 4029 2363 4063
rect 6653 4029 6687 4063
rect 10609 4029 10643 4063
rect 13277 4029 13311 4063
rect 3801 3893 3835 3927
rect 8125 3893 8159 3927
rect 12173 3689 12207 3723
rect 14657 3689 14691 3723
rect 16129 3689 16163 3723
rect 3065 3621 3099 3655
rect 5733 3621 5767 3655
rect 7941 3621 7975 3655
rect 15117 3621 15151 3655
rect 3985 3553 4019 3587
rect 10425 3553 10459 3587
rect 14749 3553 14783 3587
rect 1961 3485 1995 3519
rect 2421 3485 2455 3519
rect 6193 3485 6227 3519
rect 8953 3485 8987 3519
rect 14933 3485 14967 3519
rect 16221 3485 16255 3519
rect 4261 3417 4295 3451
rect 6469 3417 6503 3451
rect 10701 3417 10735 3451
rect 14657 3417 14691 3451
rect 1869 3349 1903 3383
rect 14473 3145 14507 3179
rect 2789 3077 2823 3111
rect 4353 3077 4387 3111
rect 8493 3077 8527 3111
rect 15117 3077 15151 3111
rect 4997 3009 5031 3043
rect 5825 3009 5859 3043
rect 6561 3009 6595 3043
rect 8217 3009 8251 3043
rect 10793 3009 10827 3043
rect 14565 3009 14599 3043
rect 15209 3009 15243 3043
rect 9965 2941 9999 2975
rect 3249 2601 3283 2635
rect 23305 2533 23339 2567
rect 1501 2465 1535 2499
rect 1777 2329 1811 2363
rect 22845 2329 22879 2363
rect 23489 2329 23523 2363
<< metal1 >>
rect 1104 27770 28888 27792
rect 1104 27718 4424 27770
rect 4476 27718 4488 27770
rect 4540 27718 4552 27770
rect 4604 27718 4616 27770
rect 4668 27718 4680 27770
rect 4732 27718 11372 27770
rect 11424 27718 11436 27770
rect 11488 27718 11500 27770
rect 11552 27718 11564 27770
rect 11616 27718 11628 27770
rect 11680 27718 18320 27770
rect 18372 27718 18384 27770
rect 18436 27718 18448 27770
rect 18500 27718 18512 27770
rect 18564 27718 18576 27770
rect 18628 27718 25268 27770
rect 25320 27718 25332 27770
rect 25384 27718 25396 27770
rect 25448 27718 25460 27770
rect 25512 27718 25524 27770
rect 25576 27718 28888 27770
rect 1104 27696 28888 27718
rect 17681 27591 17739 27597
rect 17681 27557 17693 27591
rect 17727 27588 17739 27591
rect 18046 27588 18052 27600
rect 17727 27560 18052 27588
rect 17727 27557 17739 27560
rect 17681 27551 17739 27557
rect 18046 27548 18052 27560
rect 18104 27548 18110 27600
rect 18064 27452 18092 27548
rect 18325 27455 18383 27461
rect 18325 27452 18337 27455
rect 18064 27424 18337 27452
rect 18325 27421 18337 27424
rect 18371 27421 18383 27455
rect 18325 27415 18383 27421
rect 18138 27316 18144 27328
rect 18099 27288 18144 27316
rect 18138 27276 18144 27288
rect 18196 27276 18202 27328
rect 1104 27226 28888 27248
rect 1104 27174 7898 27226
rect 7950 27174 7962 27226
rect 8014 27174 8026 27226
rect 8078 27174 8090 27226
rect 8142 27174 8154 27226
rect 8206 27174 14846 27226
rect 14898 27174 14910 27226
rect 14962 27174 14974 27226
rect 15026 27174 15038 27226
rect 15090 27174 15102 27226
rect 15154 27174 21794 27226
rect 21846 27174 21858 27226
rect 21910 27174 21922 27226
rect 21974 27174 21986 27226
rect 22038 27174 22050 27226
rect 22102 27174 28888 27226
rect 1104 27152 28888 27174
rect 1104 26682 28888 26704
rect 1104 26630 4424 26682
rect 4476 26630 4488 26682
rect 4540 26630 4552 26682
rect 4604 26630 4616 26682
rect 4668 26630 4680 26682
rect 4732 26630 11372 26682
rect 11424 26630 11436 26682
rect 11488 26630 11500 26682
rect 11552 26630 11564 26682
rect 11616 26630 11628 26682
rect 11680 26630 18320 26682
rect 18372 26630 18384 26682
rect 18436 26630 18448 26682
rect 18500 26630 18512 26682
rect 18564 26630 18576 26682
rect 18628 26630 25268 26682
rect 25320 26630 25332 26682
rect 25384 26630 25396 26682
rect 25448 26630 25460 26682
rect 25512 26630 25524 26682
rect 25576 26630 28888 26682
rect 1104 26608 28888 26630
rect 1104 26138 28888 26160
rect 1104 26086 7898 26138
rect 7950 26086 7962 26138
rect 8014 26086 8026 26138
rect 8078 26086 8090 26138
rect 8142 26086 8154 26138
rect 8206 26086 14846 26138
rect 14898 26086 14910 26138
rect 14962 26086 14974 26138
rect 15026 26086 15038 26138
rect 15090 26086 15102 26138
rect 15154 26086 21794 26138
rect 21846 26086 21858 26138
rect 21910 26086 21922 26138
rect 21974 26086 21986 26138
rect 22038 26086 22050 26138
rect 22102 26086 28888 26138
rect 1104 26064 28888 26086
rect 1104 25594 28888 25616
rect 1104 25542 4424 25594
rect 4476 25542 4488 25594
rect 4540 25542 4552 25594
rect 4604 25542 4616 25594
rect 4668 25542 4680 25594
rect 4732 25542 11372 25594
rect 11424 25542 11436 25594
rect 11488 25542 11500 25594
rect 11552 25542 11564 25594
rect 11616 25542 11628 25594
rect 11680 25542 18320 25594
rect 18372 25542 18384 25594
rect 18436 25542 18448 25594
rect 18500 25542 18512 25594
rect 18564 25542 18576 25594
rect 18628 25542 25268 25594
rect 25320 25542 25332 25594
rect 25384 25542 25396 25594
rect 25448 25542 25460 25594
rect 25512 25542 25524 25594
rect 25576 25542 28888 25594
rect 1104 25520 28888 25542
rect 1104 25050 28888 25072
rect 1104 24998 7898 25050
rect 7950 24998 7962 25050
rect 8014 24998 8026 25050
rect 8078 24998 8090 25050
rect 8142 24998 8154 25050
rect 8206 24998 14846 25050
rect 14898 24998 14910 25050
rect 14962 24998 14974 25050
rect 15026 24998 15038 25050
rect 15090 24998 15102 25050
rect 15154 24998 21794 25050
rect 21846 24998 21858 25050
rect 21910 24998 21922 25050
rect 21974 24998 21986 25050
rect 22038 24998 22050 25050
rect 22102 24998 28888 25050
rect 1104 24976 28888 24998
rect 1673 24803 1731 24809
rect 1673 24769 1685 24803
rect 1719 24800 1731 24803
rect 6362 24800 6368 24812
rect 1719 24772 6368 24800
rect 1719 24769 1731 24772
rect 1673 24763 1731 24769
rect 6362 24760 6368 24772
rect 6420 24760 6426 24812
rect 1486 24596 1492 24608
rect 1447 24568 1492 24596
rect 1486 24556 1492 24568
rect 1544 24556 1550 24608
rect 1104 24506 28888 24528
rect 1104 24454 4424 24506
rect 4476 24454 4488 24506
rect 4540 24454 4552 24506
rect 4604 24454 4616 24506
rect 4668 24454 4680 24506
rect 4732 24454 11372 24506
rect 11424 24454 11436 24506
rect 11488 24454 11500 24506
rect 11552 24454 11564 24506
rect 11616 24454 11628 24506
rect 11680 24454 18320 24506
rect 18372 24454 18384 24506
rect 18436 24454 18448 24506
rect 18500 24454 18512 24506
rect 18564 24454 18576 24506
rect 18628 24454 25268 24506
rect 25320 24454 25332 24506
rect 25384 24454 25396 24506
rect 25448 24454 25460 24506
rect 25512 24454 25524 24506
rect 25576 24454 28888 24506
rect 1104 24432 28888 24454
rect 1104 23962 28888 23984
rect 1104 23910 7898 23962
rect 7950 23910 7962 23962
rect 8014 23910 8026 23962
rect 8078 23910 8090 23962
rect 8142 23910 8154 23962
rect 8206 23910 14846 23962
rect 14898 23910 14910 23962
rect 14962 23910 14974 23962
rect 15026 23910 15038 23962
rect 15090 23910 15102 23962
rect 15154 23910 21794 23962
rect 21846 23910 21858 23962
rect 21910 23910 21922 23962
rect 21974 23910 21986 23962
rect 22038 23910 22050 23962
rect 22102 23910 28888 23962
rect 1104 23888 28888 23910
rect 1104 23418 28888 23440
rect 1104 23366 4424 23418
rect 4476 23366 4488 23418
rect 4540 23366 4552 23418
rect 4604 23366 4616 23418
rect 4668 23366 4680 23418
rect 4732 23366 11372 23418
rect 11424 23366 11436 23418
rect 11488 23366 11500 23418
rect 11552 23366 11564 23418
rect 11616 23366 11628 23418
rect 11680 23366 18320 23418
rect 18372 23366 18384 23418
rect 18436 23366 18448 23418
rect 18500 23366 18512 23418
rect 18564 23366 18576 23418
rect 18628 23366 25268 23418
rect 25320 23366 25332 23418
rect 25384 23366 25396 23418
rect 25448 23366 25460 23418
rect 25512 23366 25524 23418
rect 25576 23366 28888 23418
rect 1104 23344 28888 23366
rect 1104 22874 28888 22896
rect 1104 22822 7898 22874
rect 7950 22822 7962 22874
rect 8014 22822 8026 22874
rect 8078 22822 8090 22874
rect 8142 22822 8154 22874
rect 8206 22822 14846 22874
rect 14898 22822 14910 22874
rect 14962 22822 14974 22874
rect 15026 22822 15038 22874
rect 15090 22822 15102 22874
rect 15154 22822 21794 22874
rect 21846 22822 21858 22874
rect 21910 22822 21922 22874
rect 21974 22822 21986 22874
rect 22038 22822 22050 22874
rect 22102 22822 28888 22874
rect 1104 22800 28888 22822
rect 1104 22330 28888 22352
rect 1104 22278 4424 22330
rect 4476 22278 4488 22330
rect 4540 22278 4552 22330
rect 4604 22278 4616 22330
rect 4668 22278 4680 22330
rect 4732 22278 11372 22330
rect 11424 22278 11436 22330
rect 11488 22278 11500 22330
rect 11552 22278 11564 22330
rect 11616 22278 11628 22330
rect 11680 22278 18320 22330
rect 18372 22278 18384 22330
rect 18436 22278 18448 22330
rect 18500 22278 18512 22330
rect 18564 22278 18576 22330
rect 18628 22278 25268 22330
rect 25320 22278 25332 22330
rect 25384 22278 25396 22330
rect 25448 22278 25460 22330
rect 25512 22278 25524 22330
rect 25576 22278 28888 22330
rect 1104 22256 28888 22278
rect 1104 21786 28888 21808
rect 1104 21734 7898 21786
rect 7950 21734 7962 21786
rect 8014 21734 8026 21786
rect 8078 21734 8090 21786
rect 8142 21734 8154 21786
rect 8206 21734 14846 21786
rect 14898 21734 14910 21786
rect 14962 21734 14974 21786
rect 15026 21734 15038 21786
rect 15090 21734 15102 21786
rect 15154 21734 21794 21786
rect 21846 21734 21858 21786
rect 21910 21734 21922 21786
rect 21974 21734 21986 21786
rect 22038 21734 22050 21786
rect 22102 21734 28888 21786
rect 1104 21712 28888 21734
rect 1104 21242 28888 21264
rect 1104 21190 4424 21242
rect 4476 21190 4488 21242
rect 4540 21190 4552 21242
rect 4604 21190 4616 21242
rect 4668 21190 4680 21242
rect 4732 21190 11372 21242
rect 11424 21190 11436 21242
rect 11488 21190 11500 21242
rect 11552 21190 11564 21242
rect 11616 21190 11628 21242
rect 11680 21190 18320 21242
rect 18372 21190 18384 21242
rect 18436 21190 18448 21242
rect 18500 21190 18512 21242
rect 18564 21190 18576 21242
rect 18628 21190 25268 21242
rect 25320 21190 25332 21242
rect 25384 21190 25396 21242
rect 25448 21190 25460 21242
rect 25512 21190 25524 21242
rect 25576 21190 28888 21242
rect 1104 21168 28888 21190
rect 1104 20698 28888 20720
rect 1104 20646 7898 20698
rect 7950 20646 7962 20698
rect 8014 20646 8026 20698
rect 8078 20646 8090 20698
rect 8142 20646 8154 20698
rect 8206 20646 14846 20698
rect 14898 20646 14910 20698
rect 14962 20646 14974 20698
rect 15026 20646 15038 20698
rect 15090 20646 15102 20698
rect 15154 20646 21794 20698
rect 21846 20646 21858 20698
rect 21910 20646 21922 20698
rect 21974 20646 21986 20698
rect 22038 20646 22050 20698
rect 22102 20646 28888 20698
rect 1104 20624 28888 20646
rect 3513 20451 3571 20457
rect 3513 20417 3525 20451
rect 3559 20448 3571 20451
rect 3970 20448 3976 20460
rect 3559 20420 3976 20448
rect 3559 20417 3571 20420
rect 3513 20411 3571 20417
rect 3970 20408 3976 20420
rect 4028 20408 4034 20460
rect 3421 20247 3479 20253
rect 3421 20213 3433 20247
rect 3467 20244 3479 20247
rect 3786 20244 3792 20256
rect 3467 20216 3792 20244
rect 3467 20213 3479 20216
rect 3421 20207 3479 20213
rect 3786 20204 3792 20216
rect 3844 20204 3850 20256
rect 3970 20244 3976 20256
rect 3931 20216 3976 20244
rect 3970 20204 3976 20216
rect 4028 20204 4034 20256
rect 1104 20154 28888 20176
rect 1104 20102 4424 20154
rect 4476 20102 4488 20154
rect 4540 20102 4552 20154
rect 4604 20102 4616 20154
rect 4668 20102 4680 20154
rect 4732 20102 11372 20154
rect 11424 20102 11436 20154
rect 11488 20102 11500 20154
rect 11552 20102 11564 20154
rect 11616 20102 11628 20154
rect 11680 20102 18320 20154
rect 18372 20102 18384 20154
rect 18436 20102 18448 20154
rect 18500 20102 18512 20154
rect 18564 20102 18576 20154
rect 18628 20102 25268 20154
rect 25320 20102 25332 20154
rect 25384 20102 25396 20154
rect 25448 20102 25460 20154
rect 25512 20102 25524 20154
rect 25576 20102 28888 20154
rect 1104 20080 28888 20102
rect 2777 19839 2835 19845
rect 2777 19805 2789 19839
rect 2823 19836 2835 19839
rect 3142 19836 3148 19848
rect 2823 19808 3148 19836
rect 2823 19805 2835 19808
rect 2777 19799 2835 19805
rect 3142 19796 3148 19808
rect 3200 19836 3206 19848
rect 3789 19839 3847 19845
rect 3789 19836 3801 19839
rect 3200 19808 3801 19836
rect 3200 19796 3206 19808
rect 3789 19805 3801 19808
rect 3835 19836 3847 19839
rect 3970 19836 3976 19848
rect 3835 19808 3976 19836
rect 3835 19805 3847 19808
rect 3789 19799 3847 19805
rect 3970 19796 3976 19808
rect 4028 19796 4034 19848
rect 2869 19703 2927 19709
rect 2869 19669 2881 19703
rect 2915 19700 2927 19703
rect 3418 19700 3424 19712
rect 2915 19672 3424 19700
rect 2915 19669 2927 19672
rect 2869 19663 2927 19669
rect 3418 19660 3424 19672
rect 3476 19660 3482 19712
rect 1104 19610 28888 19632
rect 1104 19558 7898 19610
rect 7950 19558 7962 19610
rect 8014 19558 8026 19610
rect 8078 19558 8090 19610
rect 8142 19558 8154 19610
rect 8206 19558 14846 19610
rect 14898 19558 14910 19610
rect 14962 19558 14974 19610
rect 15026 19558 15038 19610
rect 15090 19558 15102 19610
rect 15154 19558 21794 19610
rect 21846 19558 21858 19610
rect 21910 19558 21922 19610
rect 21974 19558 21986 19610
rect 22038 19558 22050 19610
rect 22102 19558 28888 19610
rect 1104 19536 28888 19558
rect 1104 19066 28888 19088
rect 1104 19014 4424 19066
rect 4476 19014 4488 19066
rect 4540 19014 4552 19066
rect 4604 19014 4616 19066
rect 4668 19014 4680 19066
rect 4732 19014 11372 19066
rect 11424 19014 11436 19066
rect 11488 19014 11500 19066
rect 11552 19014 11564 19066
rect 11616 19014 11628 19066
rect 11680 19014 18320 19066
rect 18372 19014 18384 19066
rect 18436 19014 18448 19066
rect 18500 19014 18512 19066
rect 18564 19014 18576 19066
rect 18628 19014 25268 19066
rect 25320 19014 25332 19066
rect 25384 19014 25396 19066
rect 25448 19014 25460 19066
rect 25512 19014 25524 19066
rect 25576 19014 28888 19066
rect 1104 18992 28888 19014
rect 1104 18522 28888 18544
rect 1104 18470 7898 18522
rect 7950 18470 7962 18522
rect 8014 18470 8026 18522
rect 8078 18470 8090 18522
rect 8142 18470 8154 18522
rect 8206 18470 14846 18522
rect 14898 18470 14910 18522
rect 14962 18470 14974 18522
rect 15026 18470 15038 18522
rect 15090 18470 15102 18522
rect 15154 18470 21794 18522
rect 21846 18470 21858 18522
rect 21910 18470 21922 18522
rect 21974 18470 21986 18522
rect 22038 18470 22050 18522
rect 22102 18470 28888 18522
rect 1104 18448 28888 18470
rect 1104 17978 28888 18000
rect 1104 17926 4424 17978
rect 4476 17926 4488 17978
rect 4540 17926 4552 17978
rect 4604 17926 4616 17978
rect 4668 17926 4680 17978
rect 4732 17926 11372 17978
rect 11424 17926 11436 17978
rect 11488 17926 11500 17978
rect 11552 17926 11564 17978
rect 11616 17926 11628 17978
rect 11680 17926 18320 17978
rect 18372 17926 18384 17978
rect 18436 17926 18448 17978
rect 18500 17926 18512 17978
rect 18564 17926 18576 17978
rect 18628 17926 25268 17978
rect 25320 17926 25332 17978
rect 25384 17926 25396 17978
rect 25448 17926 25460 17978
rect 25512 17926 25524 17978
rect 25576 17926 28888 17978
rect 1104 17904 28888 17926
rect 1104 17434 28888 17456
rect 1104 17382 7898 17434
rect 7950 17382 7962 17434
rect 8014 17382 8026 17434
rect 8078 17382 8090 17434
rect 8142 17382 8154 17434
rect 8206 17382 14846 17434
rect 14898 17382 14910 17434
rect 14962 17382 14974 17434
rect 15026 17382 15038 17434
rect 15090 17382 15102 17434
rect 15154 17382 21794 17434
rect 21846 17382 21858 17434
rect 21910 17382 21922 17434
rect 21974 17382 21986 17434
rect 22038 17382 22050 17434
rect 22102 17382 28888 17434
rect 1104 17360 28888 17382
rect 4985 17255 5043 17261
rect 4985 17221 4997 17255
rect 5031 17252 5043 17255
rect 5626 17252 5632 17264
rect 5031 17224 5632 17252
rect 5031 17221 5043 17224
rect 4985 17215 5043 17221
rect 5626 17212 5632 17224
rect 5684 17212 5690 17264
rect 7558 17212 7564 17264
rect 7616 17252 7622 17264
rect 7616 17224 8984 17252
rect 7616 17212 7622 17224
rect 4801 17187 4859 17193
rect 4801 17153 4813 17187
rect 4847 17184 4859 17187
rect 4890 17184 4896 17196
rect 4847 17156 4896 17184
rect 4847 17153 4859 17156
rect 4801 17147 4859 17153
rect 4890 17144 4896 17156
rect 4948 17144 4954 17196
rect 8956 17193 8984 17224
rect 5077 17187 5135 17193
rect 5077 17153 5089 17187
rect 5123 17153 5135 17187
rect 5077 17147 5135 17153
rect 7837 17187 7895 17193
rect 7837 17153 7849 17187
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 8941 17187 8999 17193
rect 8941 17153 8953 17187
rect 8987 17153 8999 17187
rect 8941 17147 8999 17153
rect 27525 17187 27583 17193
rect 27525 17153 27537 17187
rect 27571 17184 27583 17187
rect 28166 17184 28172 17196
rect 27571 17156 28172 17184
rect 27571 17153 27583 17156
rect 27525 17147 27583 17153
rect 4982 17008 4988 17060
rect 5040 17048 5046 17060
rect 5092 17048 5120 17147
rect 5040 17020 5120 17048
rect 5040 17008 5046 17020
rect 7374 17008 7380 17060
rect 7432 17048 7438 17060
rect 7469 17051 7527 17057
rect 7469 17048 7481 17051
rect 7432 17020 7481 17048
rect 7432 17008 7438 17020
rect 7469 17017 7481 17020
rect 7515 17017 7527 17051
rect 7852 17048 7880 17147
rect 28166 17144 28172 17156
rect 28224 17144 28230 17196
rect 7926 17076 7932 17128
rect 7984 17116 7990 17128
rect 9030 17116 9036 17128
rect 7984 17088 8029 17116
rect 8991 17088 9036 17116
rect 7984 17076 7990 17088
rect 9030 17076 9036 17088
rect 9088 17116 9094 17128
rect 10318 17116 10324 17128
rect 9088 17088 10324 17116
rect 9088 17076 9094 17088
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 8573 17051 8631 17057
rect 8573 17048 8585 17051
rect 7852 17020 8585 17048
rect 7469 17011 7527 17017
rect 8573 17017 8585 17020
rect 8619 17017 8631 17051
rect 8573 17011 8631 17017
rect 4617 16983 4675 16989
rect 4617 16949 4629 16983
rect 4663 16980 4675 16983
rect 4798 16980 4804 16992
rect 4663 16952 4804 16980
rect 4663 16949 4675 16952
rect 4617 16943 4675 16949
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 7650 16940 7656 16992
rect 7708 16980 7714 16992
rect 10410 16980 10416 16992
rect 7708 16952 10416 16980
rect 7708 16940 7714 16952
rect 10410 16940 10416 16952
rect 10468 16940 10474 16992
rect 27982 16980 27988 16992
rect 27943 16952 27988 16980
rect 27982 16940 27988 16952
rect 28040 16940 28046 16992
rect 1104 16890 28888 16912
rect 1104 16838 4424 16890
rect 4476 16838 4488 16890
rect 4540 16838 4552 16890
rect 4604 16838 4616 16890
rect 4668 16838 4680 16890
rect 4732 16838 11372 16890
rect 11424 16838 11436 16890
rect 11488 16838 11500 16890
rect 11552 16838 11564 16890
rect 11616 16838 11628 16890
rect 11680 16838 18320 16890
rect 18372 16838 18384 16890
rect 18436 16838 18448 16890
rect 18500 16838 18512 16890
rect 18564 16838 18576 16890
rect 18628 16838 25268 16890
rect 25320 16838 25332 16890
rect 25384 16838 25396 16890
rect 25448 16838 25460 16890
rect 25512 16838 25524 16890
rect 25576 16838 28888 16890
rect 1104 16816 28888 16838
rect 7926 16736 7932 16788
rect 7984 16776 7990 16788
rect 9125 16779 9183 16785
rect 9125 16776 9137 16779
rect 7984 16748 9137 16776
rect 7984 16736 7990 16748
rect 9125 16745 9137 16748
rect 9171 16745 9183 16779
rect 9125 16739 9183 16745
rect 8220 16680 9352 16708
rect 5077 16643 5135 16649
rect 5077 16609 5089 16643
rect 5123 16640 5135 16643
rect 5626 16640 5632 16652
rect 5123 16612 5632 16640
rect 5123 16609 5135 16612
rect 5077 16603 5135 16609
rect 5626 16600 5632 16612
rect 5684 16600 5690 16652
rect 7558 16640 7564 16652
rect 7116 16612 7564 16640
rect 4798 16572 4804 16584
rect 4759 16544 4804 16572
rect 4798 16532 4804 16544
rect 4856 16532 4862 16584
rect 4982 16572 4988 16584
rect 4943 16544 4988 16572
rect 4982 16532 4988 16544
rect 5040 16532 5046 16584
rect 5169 16575 5227 16581
rect 5169 16541 5181 16575
rect 5215 16541 5227 16575
rect 5169 16535 5227 16541
rect 5353 16575 5411 16581
rect 5353 16541 5365 16575
rect 5399 16572 5411 16575
rect 5718 16572 5724 16584
rect 5399 16544 5724 16572
rect 5399 16541 5411 16544
rect 5353 16535 5411 16541
rect 2958 16464 2964 16516
rect 3016 16504 3022 16516
rect 5000 16504 5028 16532
rect 3016 16476 5028 16504
rect 5184 16504 5212 16535
rect 5718 16532 5724 16544
rect 5776 16532 5782 16584
rect 7116 16581 7144 16612
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 7742 16640 7748 16652
rect 7703 16612 7748 16640
rect 7742 16600 7748 16612
rect 7800 16600 7806 16652
rect 8220 16649 8248 16680
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16609 8263 16643
rect 8205 16603 8263 16609
rect 9324 16584 9352 16680
rect 10410 16668 10416 16720
rect 10468 16708 10474 16720
rect 10468 16680 10548 16708
rect 10468 16668 10474 16680
rect 10520 16649 10548 16680
rect 10505 16643 10563 16649
rect 9416 16612 10456 16640
rect 7101 16575 7159 16581
rect 7101 16541 7113 16575
rect 7147 16574 7159 16575
rect 8113 16575 8171 16581
rect 7147 16546 7181 16574
rect 7147 16541 7159 16546
rect 7101 16535 7159 16541
rect 8113 16541 8125 16575
rect 8159 16541 8171 16575
rect 9306 16572 9312 16584
rect 9267 16544 9312 16572
rect 8113 16535 8171 16541
rect 6638 16504 6644 16516
rect 5184 16476 6644 16504
rect 3016 16464 3022 16476
rect 4062 16396 4068 16448
rect 4120 16436 4126 16448
rect 5184 16436 5212 16476
rect 6638 16464 6644 16476
rect 6696 16464 6702 16516
rect 8128 16504 8156 16535
rect 9306 16532 9312 16544
rect 9364 16532 9370 16584
rect 9416 16581 9444 16612
rect 9401 16575 9459 16581
rect 9401 16541 9413 16575
rect 9447 16574 9459 16575
rect 9447 16546 9481 16574
rect 9582 16572 9588 16584
rect 9447 16541 9459 16546
rect 9543 16544 9588 16572
rect 9401 16535 9459 16541
rect 9416 16504 9444 16535
rect 9582 16532 9588 16544
rect 9640 16532 9646 16584
rect 9677 16575 9735 16581
rect 9677 16541 9689 16575
rect 9723 16572 9735 16575
rect 10137 16575 10195 16581
rect 10137 16572 10149 16575
rect 9723 16544 10149 16572
rect 9723 16541 9735 16544
rect 9677 16535 9735 16541
rect 10137 16541 10149 16544
rect 10183 16541 10195 16575
rect 10318 16572 10324 16584
rect 10231 16544 10324 16572
rect 10137 16535 10195 16541
rect 10318 16532 10324 16544
rect 10376 16532 10382 16584
rect 10428 16572 10456 16612
rect 10505 16609 10517 16643
rect 10551 16609 10563 16643
rect 11333 16643 11391 16649
rect 11333 16640 11345 16643
rect 10505 16603 10563 16609
rect 10612 16612 11345 16640
rect 10612 16572 10640 16612
rect 11333 16609 11345 16612
rect 11379 16609 11391 16643
rect 11333 16603 11391 16609
rect 10428 16544 10640 16572
rect 11517 16575 11575 16581
rect 11517 16541 11529 16575
rect 11563 16572 11575 16575
rect 11698 16572 11704 16584
rect 11563 16544 11704 16572
rect 11563 16541 11575 16544
rect 11517 16535 11575 16541
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 11793 16575 11851 16581
rect 11793 16541 11805 16575
rect 11839 16572 11851 16575
rect 12434 16572 12440 16584
rect 11839 16544 12440 16572
rect 11839 16541 11851 16544
rect 11793 16535 11851 16541
rect 12434 16532 12440 16544
rect 12492 16532 12498 16584
rect 10336 16504 10364 16532
rect 8128 16476 9444 16504
rect 9600 16476 10364 16504
rect 9600 16448 9628 16476
rect 5534 16436 5540 16448
rect 4120 16408 5212 16436
rect 5495 16408 5540 16436
rect 4120 16396 4126 16408
rect 5534 16396 5540 16408
rect 5592 16396 5598 16448
rect 5718 16396 5724 16448
rect 5776 16436 5782 16448
rect 7009 16439 7067 16445
rect 7009 16436 7021 16439
rect 5776 16408 7021 16436
rect 5776 16396 5782 16408
rect 7009 16405 7021 16408
rect 7055 16405 7067 16439
rect 7009 16399 7067 16405
rect 9582 16396 9588 16448
rect 9640 16396 9646 16448
rect 11698 16436 11704 16448
rect 11659 16408 11704 16436
rect 11698 16396 11704 16408
rect 11756 16396 11762 16448
rect 1104 16346 28888 16368
rect 1104 16294 7898 16346
rect 7950 16294 7962 16346
rect 8014 16294 8026 16346
rect 8078 16294 8090 16346
rect 8142 16294 8154 16346
rect 8206 16294 14846 16346
rect 14898 16294 14910 16346
rect 14962 16294 14974 16346
rect 15026 16294 15038 16346
rect 15090 16294 15102 16346
rect 15154 16294 21794 16346
rect 21846 16294 21858 16346
rect 21910 16294 21922 16346
rect 21974 16294 21986 16346
rect 22038 16294 22050 16346
rect 22102 16294 28888 16346
rect 1104 16272 28888 16294
rect 4709 16235 4767 16241
rect 4709 16201 4721 16235
rect 4755 16232 4767 16235
rect 4890 16232 4896 16244
rect 4755 16204 4896 16232
rect 4755 16201 4767 16204
rect 4709 16195 4767 16201
rect 4890 16192 4896 16204
rect 4948 16192 4954 16244
rect 7742 16192 7748 16244
rect 7800 16232 7806 16244
rect 7837 16235 7895 16241
rect 7837 16232 7849 16235
rect 7800 16204 7849 16232
rect 7800 16192 7806 16204
rect 7837 16201 7849 16204
rect 7883 16201 7895 16235
rect 9306 16232 9312 16244
rect 9267 16204 9312 16232
rect 7837 16195 7895 16201
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 5534 16124 5540 16176
rect 5592 16164 5598 16176
rect 6365 16167 6423 16173
rect 6365 16164 6377 16167
rect 5592 16136 6377 16164
rect 5592 16124 5598 16136
rect 6365 16133 6377 16136
rect 6411 16133 6423 16167
rect 6365 16127 6423 16133
rect 4890 16096 4896 16108
rect 4851 16068 4896 16096
rect 4890 16056 4896 16068
rect 4948 16056 4954 16108
rect 4982 16056 4988 16108
rect 5040 16096 5046 16108
rect 5261 16099 5319 16105
rect 5040 16068 5085 16096
rect 5040 16056 5046 16068
rect 5261 16065 5273 16099
rect 5307 16096 5319 16099
rect 5442 16096 5448 16108
rect 5307 16068 5448 16096
rect 5307 16065 5319 16068
rect 5261 16059 5319 16065
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 5718 16056 5724 16108
rect 5776 16096 5782 16108
rect 6549 16099 6607 16105
rect 6549 16096 6561 16099
rect 5776 16068 6561 16096
rect 5776 16056 5782 16068
rect 6549 16065 6561 16068
rect 6595 16065 6607 16099
rect 6549 16059 6607 16065
rect 6638 16056 6644 16108
rect 6696 16096 6702 16108
rect 6696 16068 6741 16096
rect 6696 16056 6702 16068
rect 7374 16056 7380 16108
rect 7432 16096 7438 16108
rect 8941 16099 8999 16105
rect 8941 16096 8953 16099
rect 7432 16068 8953 16096
rect 7432 16056 7438 16068
rect 8941 16065 8953 16068
rect 8987 16065 8999 16099
rect 8941 16059 8999 16065
rect 11701 16099 11759 16105
rect 11701 16065 11713 16099
rect 11747 16096 11759 16099
rect 12434 16096 12440 16108
rect 11747 16068 12440 16096
rect 11747 16065 11759 16068
rect 11701 16059 11759 16065
rect 12434 16056 12440 16068
rect 12492 16096 12498 16108
rect 12986 16096 12992 16108
rect 12492 16068 12992 16096
rect 12492 16056 12498 16068
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 3605 16031 3663 16037
rect 3605 15997 3617 16031
rect 3651 16028 3663 16031
rect 3786 16028 3792 16040
rect 3651 16000 3792 16028
rect 3651 15997 3663 16000
rect 3605 15991 3663 15997
rect 3786 15988 3792 16000
rect 3844 15988 3850 16040
rect 3881 16031 3939 16037
rect 3881 15997 3893 16031
rect 3927 16028 3939 16031
rect 4154 16028 4160 16040
rect 3927 16000 4160 16028
rect 3927 15997 3939 16000
rect 3881 15991 3939 15997
rect 4154 15988 4160 16000
rect 4212 16028 4218 16040
rect 5169 16031 5227 16037
rect 5169 16028 5181 16031
rect 4212 16000 5181 16028
rect 4212 15988 4218 16000
rect 5169 15997 5181 16000
rect 5215 15997 5227 16031
rect 5169 15991 5227 15997
rect 7466 15988 7472 16040
rect 7524 16028 7530 16040
rect 7650 16028 7656 16040
rect 7524 16000 7656 16028
rect 7524 15988 7530 16000
rect 7650 15988 7656 16000
rect 7708 16028 7714 16040
rect 7929 16031 7987 16037
rect 7929 16028 7941 16031
rect 7708 16000 7941 16028
rect 7708 15988 7714 16000
rect 7929 15997 7941 16000
rect 7975 15997 7987 16031
rect 7929 15991 7987 15997
rect 8113 16031 8171 16037
rect 8113 15997 8125 16031
rect 8159 16028 8171 16031
rect 8294 16028 8300 16040
rect 8159 16000 8300 16028
rect 8159 15997 8171 16000
rect 8113 15991 8171 15997
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 9030 16028 9036 16040
rect 8943 16000 9036 16028
rect 9030 15988 9036 16000
rect 9088 16028 9094 16040
rect 9398 16028 9404 16040
rect 9088 16000 9404 16028
rect 9088 15988 9094 16000
rect 9398 15988 9404 16000
rect 9456 15988 9462 16040
rect 6362 15960 6368 15972
rect 6323 15932 6368 15960
rect 6362 15920 6368 15932
rect 6420 15920 6426 15972
rect 7190 15852 7196 15904
rect 7248 15892 7254 15904
rect 7469 15895 7527 15901
rect 7469 15892 7481 15895
rect 7248 15864 7481 15892
rect 7248 15852 7254 15864
rect 7469 15861 7481 15864
rect 7515 15861 7527 15895
rect 11790 15892 11796 15904
rect 11751 15864 11796 15892
rect 7469 15855 7527 15861
rect 11790 15852 11796 15864
rect 11848 15852 11854 15904
rect 12158 15892 12164 15904
rect 12119 15864 12164 15892
rect 12158 15852 12164 15864
rect 12216 15852 12222 15904
rect 1104 15802 28888 15824
rect 1104 15750 4424 15802
rect 4476 15750 4488 15802
rect 4540 15750 4552 15802
rect 4604 15750 4616 15802
rect 4668 15750 4680 15802
rect 4732 15750 11372 15802
rect 11424 15750 11436 15802
rect 11488 15750 11500 15802
rect 11552 15750 11564 15802
rect 11616 15750 11628 15802
rect 11680 15750 18320 15802
rect 18372 15750 18384 15802
rect 18436 15750 18448 15802
rect 18500 15750 18512 15802
rect 18564 15750 18576 15802
rect 18628 15750 25268 15802
rect 25320 15750 25332 15802
rect 25384 15750 25396 15802
rect 25448 15750 25460 15802
rect 25512 15750 25524 15802
rect 25576 15750 28888 15802
rect 1104 15728 28888 15750
rect 5626 15648 5632 15700
rect 5684 15688 5690 15700
rect 7374 15688 7380 15700
rect 5684 15660 7380 15688
rect 5684 15648 5690 15660
rect 7374 15648 7380 15660
rect 7432 15648 7438 15700
rect 11698 15688 11704 15700
rect 9140 15660 11704 15688
rect 9140 15620 9168 15660
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 6656 15592 9168 15620
rect 9217 15623 9275 15629
rect 4982 15512 4988 15564
rect 5040 15552 5046 15564
rect 5353 15555 5411 15561
rect 5353 15552 5365 15555
rect 5040 15524 5365 15552
rect 5040 15512 5046 15524
rect 5353 15521 5365 15524
rect 5399 15552 5411 15555
rect 6549 15555 6607 15561
rect 6549 15552 6561 15555
rect 5399 15524 6561 15552
rect 5399 15521 5411 15524
rect 5353 15515 5411 15521
rect 6549 15521 6561 15524
rect 6595 15521 6607 15555
rect 6549 15515 6607 15521
rect 6656 15496 6684 15592
rect 9217 15589 9229 15623
rect 9263 15620 9275 15623
rect 9858 15620 9864 15632
rect 9263 15592 9864 15620
rect 9263 15589 9275 15592
rect 9217 15583 9275 15589
rect 9858 15580 9864 15592
rect 9916 15580 9922 15632
rect 14274 15620 14280 15632
rect 12084 15592 14280 15620
rect 6730 15512 6736 15564
rect 6788 15552 6794 15564
rect 8941 15555 8999 15561
rect 8941 15552 8953 15555
rect 6788 15524 8953 15552
rect 6788 15512 6794 15524
rect 8941 15521 8953 15524
rect 8987 15552 8999 15555
rect 9490 15552 9496 15564
rect 8987 15524 9496 15552
rect 8987 15521 8999 15524
rect 8941 15515 8999 15521
rect 9490 15512 9496 15524
rect 9548 15512 9554 15564
rect 5718 15484 5724 15496
rect 5679 15456 5724 15484
rect 5718 15444 5724 15456
rect 5776 15444 5782 15496
rect 5813 15487 5871 15493
rect 5813 15453 5825 15487
rect 5859 15484 5871 15487
rect 6362 15484 6368 15496
rect 5859 15456 6368 15484
rect 5859 15453 5871 15456
rect 5813 15447 5871 15453
rect 6362 15444 6368 15456
rect 6420 15444 6426 15496
rect 6638 15484 6644 15496
rect 6599 15456 6644 15484
rect 6638 15444 6644 15456
rect 6696 15444 6702 15496
rect 7374 15444 7380 15496
rect 7432 15484 7438 15496
rect 7469 15487 7527 15493
rect 7469 15484 7481 15487
rect 7432 15456 7481 15484
rect 7432 15444 7438 15456
rect 7469 15453 7481 15456
rect 7515 15453 7527 15487
rect 9122 15484 9128 15496
rect 9083 15456 9128 15484
rect 7469 15447 7527 15453
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 9306 15484 9312 15496
rect 9219 15456 9312 15484
rect 5997 15419 6055 15425
rect 5997 15385 6009 15419
rect 6043 15416 6055 15419
rect 9232 15416 9260 15456
rect 9306 15444 9312 15456
rect 9364 15444 9370 15496
rect 9398 15444 9404 15496
rect 9456 15484 9462 15496
rect 9456 15456 9501 15484
rect 9456 15444 9462 15456
rect 11146 15444 11152 15496
rect 11204 15484 11210 15496
rect 12084 15493 12112 15592
rect 14274 15580 14280 15592
rect 14332 15580 14338 15632
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15521 13415 15555
rect 13357 15515 13415 15521
rect 11333 15487 11391 15493
rect 11333 15484 11345 15487
rect 11204 15456 11345 15484
rect 11204 15444 11210 15456
rect 11333 15453 11345 15456
rect 11379 15484 11391 15487
rect 12069 15487 12127 15493
rect 12069 15484 12081 15487
rect 11379 15456 12081 15484
rect 11379 15453 11391 15456
rect 11333 15447 11391 15453
rect 12069 15453 12081 15456
rect 12115 15453 12127 15487
rect 12069 15447 12127 15453
rect 13372 15416 13400 15515
rect 6043 15388 9260 15416
rect 9416 15388 13400 15416
rect 6043 15385 6055 15388
rect 5997 15379 6055 15385
rect 5442 15348 5448 15360
rect 5403 15320 5448 15348
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 5626 15348 5632 15360
rect 5587 15320 5632 15348
rect 5626 15308 5632 15320
rect 5684 15308 5690 15360
rect 8294 15308 8300 15360
rect 8352 15348 8358 15360
rect 8754 15348 8760 15360
rect 8352 15320 8760 15348
rect 8352 15308 8358 15320
rect 8754 15308 8760 15320
rect 8812 15348 8818 15360
rect 9416 15348 9444 15388
rect 11882 15348 11888 15360
rect 8812 15320 9444 15348
rect 11843 15320 11888 15348
rect 8812 15308 8818 15320
rect 11882 15308 11888 15320
rect 11940 15308 11946 15360
rect 12802 15348 12808 15360
rect 12763 15320 12808 15348
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 13170 15348 13176 15360
rect 13131 15320 13176 15348
rect 13170 15308 13176 15320
rect 13228 15308 13234 15360
rect 13262 15308 13268 15360
rect 13320 15348 13326 15360
rect 13320 15320 13365 15348
rect 13320 15308 13326 15320
rect 1104 15258 28888 15280
rect 1104 15206 7898 15258
rect 7950 15206 7962 15258
rect 8014 15206 8026 15258
rect 8078 15206 8090 15258
rect 8142 15206 8154 15258
rect 8206 15206 14846 15258
rect 14898 15206 14910 15258
rect 14962 15206 14974 15258
rect 15026 15206 15038 15258
rect 15090 15206 15102 15258
rect 15154 15206 21794 15258
rect 21846 15206 21858 15258
rect 21910 15206 21922 15258
rect 21974 15206 21986 15258
rect 22038 15206 22050 15258
rect 22102 15206 28888 15258
rect 1104 15184 28888 15206
rect 4890 15144 4896 15156
rect 4851 15116 4896 15144
rect 4890 15104 4896 15116
rect 4948 15104 4954 15156
rect 5442 15104 5448 15156
rect 5500 15144 5506 15156
rect 6457 15147 6515 15153
rect 6457 15144 6469 15147
rect 5500 15116 6469 15144
rect 5500 15104 5506 15116
rect 6457 15113 6469 15116
rect 6503 15113 6515 15147
rect 6457 15107 6515 15113
rect 12621 15147 12679 15153
rect 12621 15113 12633 15147
rect 12667 15144 12679 15147
rect 13170 15144 13176 15156
rect 12667 15116 13176 15144
rect 12667 15113 12679 15116
rect 12621 15107 12679 15113
rect 13170 15104 13176 15116
rect 13228 15104 13234 15156
rect 4525 15079 4583 15085
rect 4525 15045 4537 15079
rect 4571 15076 4583 15079
rect 5460 15076 5488 15104
rect 4571 15048 5488 15076
rect 4571 15045 4583 15048
rect 4525 15039 4583 15045
rect 1946 14968 1952 15020
rect 2004 15008 2010 15020
rect 2133 15011 2191 15017
rect 2133 15008 2145 15011
rect 2004 14980 2145 15008
rect 2004 14968 2010 14980
rect 2133 14977 2145 14980
rect 2179 14977 2191 15011
rect 2133 14971 2191 14977
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 15008 2375 15011
rect 2406 15008 2412 15020
rect 2363 14980 2412 15008
rect 2363 14977 2375 14980
rect 2317 14971 2375 14977
rect 2406 14968 2412 14980
rect 2464 14968 2470 15020
rect 4154 14968 4160 15020
rect 4212 15008 4218 15020
rect 4433 15011 4491 15017
rect 4433 15008 4445 15011
rect 4212 14980 4445 15008
rect 4212 14968 4218 14980
rect 4433 14977 4445 14980
rect 4479 14977 4491 15011
rect 4433 14971 4491 14977
rect 4709 15011 4767 15017
rect 4709 14977 4721 15011
rect 4755 14977 4767 15011
rect 6546 15008 6552 15020
rect 6507 14980 6552 15008
rect 4709 14971 4767 14977
rect 3602 14900 3608 14952
rect 3660 14940 3666 14952
rect 4724 14940 4752 14971
rect 6546 14968 6552 14980
rect 6604 14968 6610 15020
rect 11698 14968 11704 15020
rect 11756 15008 11762 15020
rect 12253 15011 12311 15017
rect 12253 15008 12265 15011
rect 11756 14980 12265 15008
rect 11756 14968 11762 14980
rect 12253 14977 12265 14980
rect 12299 14977 12311 15011
rect 12253 14971 12311 14977
rect 12158 14940 12164 14952
rect 3660 14912 4752 14940
rect 12119 14912 12164 14940
rect 3660 14900 3666 14912
rect 12158 14900 12164 14912
rect 12216 14900 12222 14952
rect 2038 14764 2044 14816
rect 2096 14804 2102 14816
rect 2133 14807 2191 14813
rect 2133 14804 2145 14807
rect 2096 14776 2145 14804
rect 2096 14764 2102 14776
rect 2133 14773 2145 14776
rect 2179 14773 2191 14807
rect 7742 14804 7748 14816
rect 7655 14776 7748 14804
rect 2133 14767 2191 14773
rect 7742 14764 7748 14776
rect 7800 14804 7806 14816
rect 27982 14804 27988 14816
rect 7800 14776 27988 14804
rect 7800 14764 7806 14776
rect 27982 14764 27988 14776
rect 28040 14764 28046 14816
rect 1104 14714 28888 14736
rect 1104 14662 4424 14714
rect 4476 14662 4488 14714
rect 4540 14662 4552 14714
rect 4604 14662 4616 14714
rect 4668 14662 4680 14714
rect 4732 14662 11372 14714
rect 11424 14662 11436 14714
rect 11488 14662 11500 14714
rect 11552 14662 11564 14714
rect 11616 14662 11628 14714
rect 11680 14662 18320 14714
rect 18372 14662 18384 14714
rect 18436 14662 18448 14714
rect 18500 14662 18512 14714
rect 18564 14662 18576 14714
rect 18628 14662 25268 14714
rect 25320 14662 25332 14714
rect 25384 14662 25396 14714
rect 25448 14662 25460 14714
rect 25512 14662 25524 14714
rect 25576 14662 28888 14714
rect 1104 14640 28888 14662
rect 7377 14603 7435 14609
rect 7377 14569 7389 14603
rect 7423 14600 7435 14603
rect 9030 14600 9036 14612
rect 7423 14572 9036 14600
rect 7423 14569 7435 14572
rect 7377 14563 7435 14569
rect 2501 14535 2559 14541
rect 2501 14501 2513 14535
rect 2547 14532 2559 14535
rect 2866 14532 2872 14544
rect 2547 14504 2872 14532
rect 2547 14501 2559 14504
rect 2501 14495 2559 14501
rect 2866 14492 2872 14504
rect 2924 14532 2930 14544
rect 3786 14532 3792 14544
rect 2924 14504 3792 14532
rect 2924 14492 2930 14504
rect 3786 14492 3792 14504
rect 3844 14492 3850 14544
rect 4065 14535 4123 14541
rect 4065 14501 4077 14535
rect 4111 14501 4123 14535
rect 4065 14495 4123 14501
rect 4080 14464 4108 14495
rect 2332 14436 4108 14464
rect 2332 14405 2360 14436
rect 6546 14424 6552 14476
rect 6604 14464 6610 14476
rect 7392 14464 7420 14563
rect 9030 14560 9036 14572
rect 9088 14600 9094 14612
rect 11790 14600 11796 14612
rect 9088 14572 11192 14600
rect 11751 14572 11796 14600
rect 9088 14560 9094 14572
rect 10870 14532 10876 14544
rect 6604 14436 7420 14464
rect 8404 14504 10876 14532
rect 6604 14424 6610 14436
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14365 2375 14399
rect 2317 14359 2375 14365
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14365 2651 14399
rect 3234 14396 3240 14408
rect 3195 14368 3240 14396
rect 2593 14359 2651 14365
rect 2608 14328 2636 14359
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 3786 14396 3792 14408
rect 3747 14368 3792 14396
rect 3786 14356 3792 14368
rect 3844 14356 3850 14408
rect 4062 14396 4068 14408
rect 4023 14368 4068 14396
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 5074 14356 5080 14408
rect 5132 14396 5138 14408
rect 5169 14399 5227 14405
rect 5169 14396 5181 14399
rect 5132 14368 5181 14396
rect 5132 14356 5138 14368
rect 5169 14365 5181 14368
rect 5215 14365 5227 14399
rect 5169 14359 5227 14365
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14396 6699 14399
rect 7190 14396 7196 14408
rect 6687 14368 7196 14396
rect 6687 14365 6699 14368
rect 6641 14359 6699 14365
rect 7190 14356 7196 14368
rect 7248 14356 7254 14408
rect 7282 14356 7288 14408
rect 7340 14396 7346 14408
rect 7558 14396 7564 14408
rect 7340 14368 7385 14396
rect 7519 14368 7564 14396
rect 7340 14356 7346 14368
rect 7558 14356 7564 14368
rect 7616 14356 7622 14408
rect 8404 14405 8432 14504
rect 10870 14492 10876 14504
rect 10928 14492 10934 14544
rect 11164 14532 11192 14572
rect 11790 14560 11796 14572
rect 11848 14560 11854 14612
rect 13262 14532 13268 14544
rect 11164 14504 13268 14532
rect 8389 14399 8447 14405
rect 8389 14365 8401 14399
rect 8435 14365 8447 14399
rect 8389 14359 8447 14365
rect 9490 14356 9496 14408
rect 9548 14396 9554 14408
rect 10689 14399 10747 14405
rect 10689 14396 10701 14399
rect 9548 14368 10701 14396
rect 9548 14356 9554 14368
rect 10689 14365 10701 14368
rect 10735 14365 10747 14399
rect 10689 14359 10747 14365
rect 10781 14399 10839 14405
rect 10781 14365 10793 14399
rect 10827 14396 10839 14399
rect 10870 14396 10876 14408
rect 10827 14368 10876 14396
rect 10827 14365 10839 14368
rect 10781 14359 10839 14365
rect 10870 14356 10876 14368
rect 10928 14356 10934 14408
rect 11164 14396 11192 14504
rect 13262 14492 13268 14504
rect 13320 14492 13326 14544
rect 11514 14464 11520 14476
rect 11475 14436 11520 14464
rect 11514 14424 11520 14436
rect 11572 14424 11578 14476
rect 11333 14399 11391 14405
rect 11333 14396 11345 14399
rect 11164 14368 11345 14396
rect 11333 14365 11345 14368
rect 11379 14365 11391 14399
rect 11333 14359 11391 14365
rect 11422 14356 11428 14408
rect 11480 14396 11486 14408
rect 11609 14399 11667 14405
rect 11480 14368 11525 14396
rect 11480 14356 11486 14368
rect 11609 14365 11621 14399
rect 11655 14365 11667 14399
rect 11609 14359 11667 14365
rect 12437 14399 12495 14405
rect 12437 14365 12449 14399
rect 12483 14396 12495 14399
rect 12526 14396 12532 14408
rect 12483 14368 12532 14396
rect 12483 14365 12495 14368
rect 12437 14359 12495 14365
rect 2682 14328 2688 14340
rect 2595 14300 2688 14328
rect 2682 14288 2688 14300
rect 2740 14328 2746 14340
rect 8297 14331 8355 14337
rect 8297 14328 8309 14331
rect 2740 14300 3924 14328
rect 2740 14288 2746 14300
rect 3896 14272 3924 14300
rect 7300 14300 8309 14328
rect 7300 14272 7328 14300
rect 8297 14297 8309 14300
rect 8343 14297 8355 14331
rect 9858 14328 9864 14340
rect 9819 14300 9864 14328
rect 8297 14291 8355 14297
rect 9858 14288 9864 14300
rect 9916 14288 9922 14340
rect 11054 14288 11060 14340
rect 11112 14328 11118 14340
rect 11624 14328 11652 14359
rect 12526 14356 12532 14368
rect 12584 14356 12590 14408
rect 12342 14328 12348 14340
rect 11112 14300 12348 14328
rect 11112 14288 11118 14300
rect 12342 14288 12348 14300
rect 12400 14288 12406 14340
rect 2130 14260 2136 14272
rect 2091 14232 2136 14260
rect 2130 14220 2136 14232
rect 2188 14220 2194 14272
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 3053 14263 3111 14269
rect 3053 14260 3065 14263
rect 2832 14232 3065 14260
rect 2832 14220 2838 14232
rect 3053 14229 3065 14232
rect 3099 14229 3111 14263
rect 3878 14260 3884 14272
rect 3839 14232 3884 14260
rect 3053 14223 3111 14229
rect 3878 14220 3884 14232
rect 3936 14220 3942 14272
rect 3970 14220 3976 14272
rect 4028 14260 4034 14272
rect 5077 14263 5135 14269
rect 5077 14260 5089 14263
rect 4028 14232 5089 14260
rect 4028 14220 4034 14232
rect 5077 14229 5089 14232
rect 5123 14229 5135 14263
rect 6454 14260 6460 14272
rect 6415 14232 6460 14260
rect 5077 14223 5135 14229
rect 6454 14220 6460 14232
rect 6512 14220 6518 14272
rect 7282 14220 7288 14272
rect 7340 14220 7346 14272
rect 7745 14263 7803 14269
rect 7745 14229 7757 14263
rect 7791 14260 7803 14263
rect 9674 14260 9680 14272
rect 7791 14232 9680 14260
rect 7791 14229 7803 14232
rect 7745 14223 7803 14229
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 9769 14263 9827 14269
rect 9769 14229 9781 14263
rect 9815 14260 9827 14263
rect 10042 14260 10048 14272
rect 9815 14232 10048 14260
rect 9815 14229 9827 14232
rect 9769 14223 9827 14229
rect 10042 14220 10048 14232
rect 10100 14260 10106 14272
rect 12250 14260 12256 14272
rect 10100 14232 12256 14260
rect 10100 14220 10106 14232
rect 12250 14220 12256 14232
rect 12308 14220 12314 14272
rect 1104 14170 28888 14192
rect 1104 14118 7898 14170
rect 7950 14118 7962 14170
rect 8014 14118 8026 14170
rect 8078 14118 8090 14170
rect 8142 14118 8154 14170
rect 8206 14118 14846 14170
rect 14898 14118 14910 14170
rect 14962 14118 14974 14170
rect 15026 14118 15038 14170
rect 15090 14118 15102 14170
rect 15154 14118 21794 14170
rect 21846 14118 21858 14170
rect 21910 14118 21922 14170
rect 21974 14118 21986 14170
rect 22038 14118 22050 14170
rect 22102 14118 28888 14170
rect 1104 14096 28888 14118
rect 2133 14059 2191 14065
rect 2133 14025 2145 14059
rect 2179 14056 2191 14059
rect 3234 14056 3240 14068
rect 2179 14028 3240 14056
rect 2179 14025 2191 14028
rect 2133 14019 2191 14025
rect 3234 14016 3240 14028
rect 3292 14016 3298 14068
rect 7193 14059 7251 14065
rect 7193 14025 7205 14059
rect 7239 14056 7251 14059
rect 7742 14056 7748 14068
rect 7239 14028 7748 14056
rect 7239 14025 7251 14028
rect 7193 14019 7251 14025
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 8754 14056 8760 14068
rect 8715 14028 8760 14056
rect 8754 14016 8760 14028
rect 8812 14016 8818 14068
rect 9582 14016 9588 14068
rect 9640 14056 9646 14068
rect 10321 14059 10379 14065
rect 10321 14056 10333 14059
rect 9640 14028 10333 14056
rect 9640 14016 9646 14028
rect 10321 14025 10333 14028
rect 10367 14025 10379 14059
rect 12986 14056 12992 14068
rect 12947 14028 12992 14056
rect 10321 14019 10379 14025
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 3142 13988 3148 14000
rect 3055 13960 3148 13988
rect 2777 13923 2835 13929
rect 2777 13889 2789 13923
rect 2823 13889 2835 13923
rect 2777 13883 2835 13889
rect 1670 13852 1676 13864
rect 1583 13824 1676 13852
rect 1670 13812 1676 13824
rect 1728 13852 1734 13864
rect 2593 13855 2651 13861
rect 2593 13852 2605 13855
rect 1728 13824 2605 13852
rect 1728 13812 1734 13824
rect 2593 13821 2605 13824
rect 2639 13821 2651 13855
rect 2792 13852 2820 13883
rect 2866 13880 2872 13932
rect 2924 13920 2930 13932
rect 3068 13929 3096 13960
rect 3142 13948 3148 13960
rect 3200 13988 3206 14000
rect 4062 13988 4068 14000
rect 3200 13960 4068 13988
rect 3200 13948 3206 13960
rect 4062 13948 4068 13960
rect 4120 13948 4126 14000
rect 6638 13988 6644 14000
rect 5460 13960 6644 13988
rect 3053 13923 3111 13929
rect 2924 13892 2969 13920
rect 2924 13880 2930 13892
rect 3053 13889 3065 13923
rect 3099 13889 3111 13923
rect 3878 13920 3884 13932
rect 3839 13892 3884 13920
rect 3053 13883 3111 13889
rect 3878 13880 3884 13892
rect 3936 13880 3942 13932
rect 5460 13929 5488 13960
rect 6638 13948 6644 13960
rect 6696 13948 6702 14000
rect 9674 13948 9680 14000
rect 9732 13988 9738 14000
rect 9861 13991 9919 13997
rect 9861 13988 9873 13991
rect 9732 13960 9873 13988
rect 9732 13948 9738 13960
rect 9861 13957 9873 13960
rect 9907 13957 9919 13991
rect 9861 13951 9919 13957
rect 11422 13948 11428 14000
rect 11480 13988 11486 14000
rect 13449 13991 13507 13997
rect 13449 13988 13461 13991
rect 11480 13960 13461 13988
rect 11480 13948 11486 13960
rect 13449 13957 13461 13960
rect 13495 13957 13507 13991
rect 13449 13951 13507 13957
rect 5445 13923 5503 13929
rect 5445 13889 5457 13923
rect 5491 13889 5503 13923
rect 5445 13883 5503 13889
rect 6546 13880 6552 13932
rect 6604 13920 6610 13932
rect 8021 13923 8079 13929
rect 6604 13892 7144 13920
rect 6604 13880 6610 13892
rect 3234 13852 3240 13864
rect 2792 13824 3240 13852
rect 2593 13815 2651 13821
rect 3234 13812 3240 13824
rect 3292 13852 3298 13864
rect 3602 13852 3608 13864
rect 3292 13824 3608 13852
rect 3292 13812 3298 13824
rect 3602 13812 3608 13824
rect 3660 13812 3666 13864
rect 5353 13855 5411 13861
rect 5353 13821 5365 13855
rect 5399 13852 5411 13855
rect 6730 13852 6736 13864
rect 5399 13824 6736 13852
rect 5399 13821 5411 13824
rect 5353 13815 5411 13821
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 7116 13861 7144 13892
rect 8021 13889 8033 13923
rect 8067 13889 8079 13923
rect 8021 13883 8079 13889
rect 8113 13923 8171 13929
rect 8113 13889 8125 13923
rect 8159 13920 8171 13923
rect 8941 13923 8999 13929
rect 8941 13920 8953 13923
rect 8159 13892 8953 13920
rect 8159 13889 8171 13892
rect 8113 13883 8171 13889
rect 8941 13889 8953 13892
rect 8987 13920 8999 13923
rect 9122 13920 9128 13932
rect 8987 13892 9128 13920
rect 8987 13889 8999 13892
rect 8941 13883 8999 13889
rect 7009 13855 7067 13861
rect 7009 13821 7021 13855
rect 7055 13821 7067 13855
rect 7009 13815 7067 13821
rect 7101 13855 7159 13861
rect 7101 13821 7113 13855
rect 7147 13852 7159 13855
rect 8036 13852 8064 13883
rect 9122 13880 9128 13892
rect 9180 13880 9186 13932
rect 9217 13923 9275 13929
rect 9217 13889 9229 13923
rect 9263 13920 9275 13923
rect 9766 13920 9772 13932
rect 9263 13892 9772 13920
rect 9263 13889 9275 13892
rect 9217 13883 9275 13889
rect 9766 13880 9772 13892
rect 9824 13880 9830 13932
rect 10137 13923 10195 13929
rect 10137 13920 10149 13923
rect 9876 13892 10149 13920
rect 9876 13864 9904 13892
rect 10137 13889 10149 13892
rect 10183 13889 10195 13923
rect 10137 13883 10195 13889
rect 12342 13880 12348 13932
rect 12400 13920 12406 13932
rect 13173 13923 13231 13929
rect 13173 13920 13185 13923
rect 12400 13892 13185 13920
rect 12400 13880 12406 13892
rect 13173 13889 13185 13892
rect 13219 13889 13231 13923
rect 13173 13883 13231 13889
rect 13722 13880 13728 13932
rect 13780 13920 13786 13932
rect 14001 13923 14059 13929
rect 14001 13920 14013 13923
rect 13780 13892 14013 13920
rect 13780 13880 13786 13892
rect 14001 13889 14013 13892
rect 14047 13889 14059 13923
rect 14001 13883 14059 13889
rect 14093 13923 14151 13929
rect 14093 13889 14105 13923
rect 14139 13889 14151 13923
rect 14093 13883 14151 13889
rect 9306 13852 9312 13864
rect 7147 13824 8064 13852
rect 9140 13824 9312 13852
rect 7147 13821 7159 13824
rect 7101 13815 7159 13821
rect 1946 13784 1952 13796
rect 1907 13756 1952 13784
rect 1946 13744 1952 13756
rect 2004 13744 2010 13796
rect 2958 13784 2964 13796
rect 2919 13756 2964 13784
rect 2958 13744 2964 13756
rect 3016 13744 3022 13796
rect 5810 13784 5816 13796
rect 5771 13756 5816 13784
rect 5810 13744 5816 13756
rect 5868 13744 5874 13796
rect 6822 13744 6828 13796
rect 6880 13784 6886 13796
rect 7024 13784 7052 13815
rect 9140 13793 9168 13824
rect 9306 13812 9312 13824
rect 9364 13812 9370 13864
rect 9858 13812 9864 13864
rect 9916 13812 9922 13864
rect 9950 13812 9956 13864
rect 10008 13852 10014 13864
rect 11514 13852 11520 13864
rect 10008 13824 11520 13852
rect 10008 13812 10014 13824
rect 11514 13812 11520 13824
rect 11572 13852 11578 13864
rect 12253 13855 12311 13861
rect 12253 13852 12265 13855
rect 11572 13824 12265 13852
rect 11572 13812 11578 13824
rect 12253 13821 12265 13824
rect 12299 13821 12311 13855
rect 12253 13815 12311 13821
rect 12529 13855 12587 13861
rect 12529 13821 12541 13855
rect 12575 13852 12587 13855
rect 13357 13855 13415 13861
rect 13357 13852 13369 13855
rect 12575 13824 13369 13852
rect 12575 13821 12587 13824
rect 12529 13815 12587 13821
rect 13357 13821 13369 13824
rect 13403 13852 13415 13855
rect 13814 13852 13820 13864
rect 13403 13824 13820 13852
rect 13403 13821 13415 13824
rect 13357 13815 13415 13821
rect 13814 13812 13820 13824
rect 13872 13812 13878 13864
rect 14108 13796 14136 13883
rect 9033 13787 9091 13793
rect 9033 13784 9045 13787
rect 6880 13756 9045 13784
rect 6880 13744 6886 13756
rect 9033 13753 9045 13756
rect 9079 13753 9091 13787
rect 9033 13747 9091 13753
rect 9125 13787 9183 13793
rect 9125 13753 9137 13787
rect 9171 13753 9183 13787
rect 9125 13747 9183 13753
rect 7466 13676 7472 13728
rect 7524 13716 7530 13728
rect 7561 13719 7619 13725
rect 7561 13716 7573 13719
rect 7524 13688 7573 13716
rect 7524 13676 7530 13688
rect 7561 13685 7573 13688
rect 7607 13685 7619 13719
rect 9048 13716 9076 13747
rect 9398 13744 9404 13796
rect 9456 13784 9462 13796
rect 11882 13784 11888 13796
rect 9456 13756 11888 13784
rect 9456 13744 9462 13756
rect 11882 13744 11888 13756
rect 11940 13784 11946 13796
rect 14090 13784 14096 13796
rect 11940 13756 14096 13784
rect 11940 13744 11946 13756
rect 14090 13744 14096 13756
rect 14148 13744 14154 13796
rect 10042 13716 10048 13728
rect 9048 13688 10048 13716
rect 7561 13679 7619 13685
rect 10042 13676 10048 13688
rect 10100 13676 10106 13728
rect 10137 13719 10195 13725
rect 10137 13685 10149 13719
rect 10183 13716 10195 13719
rect 11054 13716 11060 13728
rect 10183 13688 11060 13716
rect 10183 13685 10195 13688
rect 10137 13679 10195 13685
rect 11054 13676 11060 13688
rect 11112 13676 11118 13728
rect 13262 13716 13268 13728
rect 13223 13688 13268 13716
rect 13262 13676 13268 13688
rect 13320 13676 13326 13728
rect 1104 13626 28888 13648
rect 1104 13574 4424 13626
rect 4476 13574 4488 13626
rect 4540 13574 4552 13626
rect 4604 13574 4616 13626
rect 4668 13574 4680 13626
rect 4732 13574 11372 13626
rect 11424 13574 11436 13626
rect 11488 13574 11500 13626
rect 11552 13574 11564 13626
rect 11616 13574 11628 13626
rect 11680 13574 18320 13626
rect 18372 13574 18384 13626
rect 18436 13574 18448 13626
rect 18500 13574 18512 13626
rect 18564 13574 18576 13626
rect 18628 13574 25268 13626
rect 25320 13574 25332 13626
rect 25384 13574 25396 13626
rect 25448 13574 25460 13626
rect 25512 13574 25524 13626
rect 25576 13574 28888 13626
rect 1104 13552 28888 13574
rect 1946 13472 1952 13524
rect 2004 13512 2010 13524
rect 2317 13515 2375 13521
rect 2317 13512 2329 13515
rect 2004 13484 2329 13512
rect 2004 13472 2010 13484
rect 2317 13481 2329 13484
rect 2363 13481 2375 13515
rect 2317 13475 2375 13481
rect 9766 13472 9772 13524
rect 9824 13512 9830 13524
rect 10505 13515 10563 13521
rect 10505 13512 10517 13515
rect 9824 13484 10517 13512
rect 9824 13472 9830 13484
rect 10505 13481 10517 13484
rect 10551 13481 10563 13515
rect 10505 13475 10563 13481
rect 10689 13515 10747 13521
rect 10689 13481 10701 13515
rect 10735 13481 10747 13515
rect 10689 13475 10747 13481
rect 9950 13404 9956 13456
rect 10008 13444 10014 13456
rect 10704 13444 10732 13475
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 14093 13515 14151 13521
rect 14093 13512 14105 13515
rect 13872 13484 14105 13512
rect 13872 13472 13878 13484
rect 14093 13481 14105 13484
rect 14139 13481 14151 13515
rect 14093 13475 14151 13481
rect 14461 13515 14519 13521
rect 14461 13481 14473 13515
rect 14507 13512 14519 13515
rect 15562 13512 15568 13524
rect 14507 13484 15568 13512
rect 14507 13481 14519 13484
rect 14461 13475 14519 13481
rect 15562 13472 15568 13484
rect 15620 13472 15626 13524
rect 10008 13416 10732 13444
rect 10008 13404 10014 13416
rect 10870 13404 10876 13456
rect 10928 13444 10934 13456
rect 15013 13447 15071 13453
rect 15013 13444 15025 13447
rect 10928 13416 15025 13444
rect 10928 13404 10934 13416
rect 15013 13413 15025 13416
rect 15059 13413 15071 13447
rect 15013 13407 15071 13413
rect 2682 13376 2688 13388
rect 1872 13348 2688 13376
rect 1670 13308 1676 13320
rect 1631 13280 1676 13308
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 1872 13317 1900 13348
rect 2682 13336 2688 13348
rect 2740 13336 2746 13388
rect 2777 13379 2835 13385
rect 2777 13345 2789 13379
rect 2823 13376 2835 13379
rect 3142 13376 3148 13388
rect 2823 13348 3148 13376
rect 2823 13345 2835 13348
rect 2777 13339 2835 13345
rect 3142 13336 3148 13348
rect 3200 13336 3206 13388
rect 6362 13336 6368 13388
rect 6420 13376 6426 13388
rect 6641 13379 6699 13385
rect 6641 13376 6653 13379
rect 6420 13348 6653 13376
rect 6420 13336 6426 13348
rect 6641 13345 6653 13348
rect 6687 13345 6699 13379
rect 6822 13376 6828 13388
rect 6783 13348 6828 13376
rect 6641 13339 6699 13345
rect 6822 13336 6828 13348
rect 6880 13336 6886 13388
rect 9766 13376 9772 13388
rect 7944 13348 9772 13376
rect 1857 13311 1915 13317
rect 1857 13277 1869 13311
rect 1903 13277 1915 13311
rect 1857 13271 1915 13277
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13277 2559 13311
rect 2501 13271 2559 13277
rect 2593 13311 2651 13317
rect 2593 13277 2605 13311
rect 2639 13277 2651 13311
rect 2593 13271 2651 13277
rect 4433 13311 4491 13317
rect 4433 13277 4445 13311
rect 4479 13308 4491 13311
rect 5074 13308 5080 13320
rect 4479 13280 5080 13308
rect 4479 13277 4491 13280
rect 4433 13271 4491 13277
rect 1762 13172 1768 13184
rect 1723 13144 1768 13172
rect 1762 13132 1768 13144
rect 1820 13132 1826 13184
rect 2516 13172 2544 13271
rect 2608 13240 2636 13271
rect 5074 13268 5080 13280
rect 5132 13268 5138 13320
rect 7944 13317 7972 13348
rect 9766 13336 9772 13348
rect 9824 13336 9830 13388
rect 10781 13379 10839 13385
rect 10781 13345 10793 13379
rect 10827 13376 10839 13379
rect 11054 13376 11060 13388
rect 10827 13348 11060 13376
rect 10827 13345 10839 13348
rect 10781 13339 10839 13345
rect 11054 13336 11060 13348
rect 11112 13336 11118 13388
rect 12342 13336 12348 13388
rect 12400 13376 12406 13388
rect 12529 13379 12587 13385
rect 12529 13376 12541 13379
rect 12400 13348 12541 13376
rect 12400 13336 12406 13348
rect 12529 13345 12541 13348
rect 12575 13345 12587 13379
rect 12529 13339 12587 13345
rect 5721 13311 5779 13317
rect 5721 13277 5733 13311
rect 5767 13308 5779 13311
rect 7929 13311 7987 13317
rect 5767 13280 6914 13308
rect 5767 13277 5779 13280
rect 5721 13271 5779 13277
rect 2866 13240 2872 13252
rect 2608 13212 2872 13240
rect 2866 13200 2872 13212
rect 2924 13200 2930 13252
rect 4246 13240 4252 13252
rect 4207 13212 4252 13240
rect 4246 13200 4252 13212
rect 4304 13200 4310 13252
rect 6886 13240 6914 13280
rect 7929 13277 7941 13311
rect 7975 13277 7987 13311
rect 7929 13271 7987 13277
rect 9033 13311 9091 13317
rect 9033 13277 9045 13311
rect 9079 13308 9091 13311
rect 9398 13308 9404 13320
rect 9079 13280 9404 13308
rect 9079 13277 9091 13280
rect 9033 13271 9091 13277
rect 9048 13240 9076 13271
rect 9398 13268 9404 13280
rect 9456 13268 9462 13320
rect 9674 13308 9680 13320
rect 9635 13280 9680 13308
rect 9674 13268 9680 13280
rect 9732 13268 9738 13320
rect 10045 13311 10103 13317
rect 10045 13277 10057 13311
rect 10091 13308 10103 13311
rect 10873 13311 10931 13317
rect 10873 13308 10885 13311
rect 10091 13280 10885 13308
rect 10091 13277 10103 13280
rect 10045 13271 10103 13277
rect 10873 13277 10885 13280
rect 10919 13308 10931 13311
rect 11238 13308 11244 13320
rect 10919 13280 11244 13308
rect 10919 13277 10931 13280
rect 10873 13271 10931 13277
rect 11238 13268 11244 13280
rect 11296 13268 11302 13320
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13308 11575 13311
rect 12802 13308 12808 13320
rect 11563 13280 12808 13308
rect 11563 13277 11575 13280
rect 11517 13271 11575 13277
rect 12802 13268 12808 13280
rect 12860 13268 12866 13320
rect 14366 13308 14372 13320
rect 14327 13280 14372 13308
rect 14366 13268 14372 13280
rect 14424 13268 14430 13320
rect 14461 13311 14519 13317
rect 14461 13277 14473 13311
rect 14507 13277 14519 13311
rect 14461 13271 14519 13277
rect 15197 13311 15255 13317
rect 15197 13277 15209 13311
rect 15243 13308 15255 13311
rect 15286 13308 15292 13320
rect 15243 13280 15292 13308
rect 15243 13277 15255 13280
rect 15197 13271 15255 13277
rect 9858 13240 9864 13252
rect 6886 13212 9076 13240
rect 9819 13212 9864 13240
rect 9858 13200 9864 13212
rect 9916 13240 9922 13252
rect 12437 13243 12495 13249
rect 12437 13240 12449 13243
rect 9916 13212 12449 13240
rect 9916 13200 9922 13212
rect 12437 13209 12449 13212
rect 12483 13209 12495 13243
rect 12437 13203 12495 13209
rect 14182 13200 14188 13252
rect 14240 13240 14246 13252
rect 14476 13240 14504 13271
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 14240 13212 14504 13240
rect 14240 13200 14246 13212
rect 2958 13172 2964 13184
rect 2516 13144 2964 13172
rect 2958 13132 2964 13144
rect 3016 13132 3022 13184
rect 4982 13172 4988 13184
rect 4943 13144 4988 13172
rect 4982 13132 4988 13144
rect 5040 13132 5046 13184
rect 5442 13132 5448 13184
rect 5500 13172 5506 13184
rect 5629 13175 5687 13181
rect 5629 13172 5641 13175
rect 5500 13144 5641 13172
rect 5500 13132 5506 13144
rect 5629 13141 5641 13144
rect 5675 13141 5687 13175
rect 6178 13172 6184 13184
rect 6139 13144 6184 13172
rect 5629 13135 5687 13141
rect 6178 13132 6184 13144
rect 6236 13132 6242 13184
rect 6546 13172 6552 13184
rect 6507 13144 6552 13172
rect 6546 13132 6552 13144
rect 6604 13132 6610 13184
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 7837 13175 7895 13181
rect 7837 13172 7849 13175
rect 7708 13144 7849 13172
rect 7708 13132 7714 13144
rect 7837 13141 7849 13144
rect 7883 13141 7895 13175
rect 7837 13135 7895 13141
rect 9125 13175 9183 13181
rect 9125 13141 9137 13175
rect 9171 13172 9183 13175
rect 10686 13172 10692 13184
rect 9171 13144 10692 13172
rect 9171 13141 9183 13144
rect 9125 13135 9183 13141
rect 10686 13132 10692 13144
rect 10744 13132 10750 13184
rect 10778 13132 10784 13184
rect 10836 13172 10842 13184
rect 11333 13175 11391 13181
rect 11333 13172 11345 13175
rect 10836 13144 11345 13172
rect 10836 13132 10842 13144
rect 11333 13141 11345 13144
rect 11379 13141 11391 13175
rect 11974 13172 11980 13184
rect 11935 13144 11980 13172
rect 11333 13135 11391 13141
rect 11974 13132 11980 13144
rect 12032 13132 12038 13184
rect 12345 13175 12403 13181
rect 12345 13141 12357 13175
rect 12391 13172 12403 13175
rect 12526 13172 12532 13184
rect 12391 13144 12532 13172
rect 12391 13141 12403 13144
rect 12345 13135 12403 13141
rect 12526 13132 12532 13144
rect 12584 13132 12590 13184
rect 1104 13082 28888 13104
rect 1104 13030 7898 13082
rect 7950 13030 7962 13082
rect 8014 13030 8026 13082
rect 8078 13030 8090 13082
rect 8142 13030 8154 13082
rect 8206 13030 14846 13082
rect 14898 13030 14910 13082
rect 14962 13030 14974 13082
rect 15026 13030 15038 13082
rect 15090 13030 15102 13082
rect 15154 13030 21794 13082
rect 21846 13030 21858 13082
rect 21910 13030 21922 13082
rect 21974 13030 21986 13082
rect 22038 13030 22050 13082
rect 22102 13030 28888 13082
rect 1104 13008 28888 13030
rect 2225 12971 2283 12977
rect 2225 12937 2237 12971
rect 2271 12968 2283 12971
rect 2682 12968 2688 12980
rect 2271 12940 2688 12968
rect 2271 12937 2283 12940
rect 2225 12931 2283 12937
rect 2682 12928 2688 12940
rect 2740 12928 2746 12980
rect 3697 12971 3755 12977
rect 3697 12937 3709 12971
rect 3743 12968 3755 12971
rect 4246 12968 4252 12980
rect 3743 12940 4252 12968
rect 3743 12937 3755 12940
rect 3697 12931 3755 12937
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 14366 12928 14372 12980
rect 14424 12968 14430 12980
rect 14737 12971 14795 12977
rect 14737 12968 14749 12971
rect 14424 12940 14749 12968
rect 14424 12928 14430 12940
rect 14737 12937 14749 12940
rect 14783 12937 14795 12971
rect 14737 12931 14795 12937
rect 2866 12900 2872 12912
rect 2148 12872 2872 12900
rect 2148 12841 2176 12872
rect 2866 12860 2872 12872
rect 2924 12860 2930 12912
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12801 2191 12835
rect 2133 12795 2191 12801
rect 2409 12835 2467 12841
rect 2409 12801 2421 12835
rect 2455 12832 2467 12835
rect 2958 12832 2964 12844
rect 2455 12804 2964 12832
rect 2455 12801 2467 12804
rect 2409 12795 2467 12801
rect 2958 12792 2964 12804
rect 3016 12832 3022 12844
rect 3326 12832 3332 12844
rect 3016 12804 3332 12832
rect 3016 12792 3022 12804
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 4341 12835 4399 12841
rect 4341 12801 4353 12835
rect 4387 12832 4399 12835
rect 4985 12835 5043 12841
rect 4985 12832 4997 12835
rect 4387 12804 4997 12832
rect 4387 12801 4399 12804
rect 4341 12795 4399 12801
rect 4985 12801 4997 12804
rect 5031 12832 5043 12835
rect 5074 12832 5080 12844
rect 5031 12804 5080 12832
rect 5031 12801 5043 12804
rect 4985 12795 5043 12801
rect 5074 12792 5080 12804
rect 5132 12832 5138 12844
rect 5445 12835 5503 12841
rect 5445 12832 5457 12835
rect 5132 12804 5457 12832
rect 5132 12792 5138 12804
rect 5445 12801 5457 12804
rect 5491 12801 5503 12835
rect 5445 12795 5503 12801
rect 7009 12835 7067 12841
rect 7009 12801 7021 12835
rect 7055 12801 7067 12835
rect 7466 12832 7472 12844
rect 7427 12804 7472 12832
rect 7009 12795 7067 12801
rect 3510 12724 3516 12776
rect 3568 12764 3574 12776
rect 4893 12767 4951 12773
rect 4893 12764 4905 12767
rect 3568 12736 4905 12764
rect 3568 12724 3574 12736
rect 4893 12733 4905 12736
rect 4939 12733 4951 12767
rect 7024 12764 7052 12795
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12832 9459 12835
rect 9766 12832 9772 12844
rect 9447 12804 9772 12832
rect 9447 12801 9459 12804
rect 9401 12795 9459 12801
rect 9416 12764 9444 12795
rect 9766 12792 9772 12804
rect 9824 12832 9830 12844
rect 10870 12832 10876 12844
rect 9824 12804 10876 12832
rect 9824 12792 9830 12804
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 11974 12832 11980 12844
rect 11935 12804 11980 12832
rect 11974 12792 11980 12804
rect 12032 12792 12038 12844
rect 14093 12835 14151 12841
rect 14093 12801 14105 12835
rect 14139 12832 14151 12835
rect 14182 12832 14188 12844
rect 14139 12804 14188 12832
rect 14139 12801 14151 12804
rect 14093 12795 14151 12801
rect 14182 12792 14188 12804
rect 14240 12792 14246 12844
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12801 14611 12835
rect 14553 12795 14611 12801
rect 7024 12736 9444 12764
rect 4893 12727 4951 12733
rect 13630 12724 13636 12776
rect 13688 12764 13694 12776
rect 13817 12767 13875 12773
rect 13817 12764 13829 12767
rect 13688 12736 13829 12764
rect 13688 12724 13694 12736
rect 13817 12733 13829 12736
rect 13863 12764 13875 12767
rect 14568 12764 14596 12795
rect 13863 12736 14596 12764
rect 13863 12733 13875 12736
rect 13817 12727 13875 12733
rect 2406 12696 2412 12708
rect 2367 12668 2412 12696
rect 2406 12656 2412 12668
rect 2464 12656 2470 12708
rect 3878 12656 3884 12708
rect 3936 12696 3942 12708
rect 5537 12699 5595 12705
rect 5537 12696 5549 12699
rect 3936 12668 5549 12696
rect 3936 12656 3942 12668
rect 5537 12665 5549 12668
rect 5583 12665 5595 12699
rect 5537 12659 5595 12665
rect 14001 12699 14059 12705
rect 14001 12665 14013 12699
rect 14047 12696 14059 12699
rect 15562 12696 15568 12708
rect 14047 12668 15568 12696
rect 14047 12665 14059 12668
rect 14001 12659 14059 12665
rect 15562 12656 15568 12668
rect 15620 12656 15626 12708
rect 4249 12631 4307 12637
rect 4249 12597 4261 12631
rect 4295 12628 4307 12631
rect 4798 12628 4804 12640
rect 4295 12600 4804 12628
rect 4295 12597 4307 12600
rect 4249 12591 4307 12597
rect 4798 12588 4804 12600
rect 4856 12588 4862 12640
rect 6914 12588 6920 12640
rect 6972 12628 6978 12640
rect 7653 12631 7711 12637
rect 6972 12600 7017 12628
rect 6972 12588 6978 12600
rect 7653 12597 7665 12631
rect 7699 12628 7711 12631
rect 7742 12628 7748 12640
rect 7699 12600 7748 12628
rect 7699 12597 7711 12600
rect 7653 12591 7711 12597
rect 7742 12588 7748 12600
rect 7800 12588 7806 12640
rect 9493 12631 9551 12637
rect 9493 12597 9505 12631
rect 9539 12628 9551 12631
rect 9674 12628 9680 12640
rect 9539 12600 9680 12628
rect 9539 12597 9551 12600
rect 9493 12591 9551 12597
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 11790 12628 11796 12640
rect 11751 12600 11796 12628
rect 11790 12588 11796 12600
rect 11848 12588 11854 12640
rect 13906 12628 13912 12640
rect 13867 12600 13912 12628
rect 13906 12588 13912 12600
rect 13964 12588 13970 12640
rect 1104 12538 28888 12560
rect 1104 12486 4424 12538
rect 4476 12486 4488 12538
rect 4540 12486 4552 12538
rect 4604 12486 4616 12538
rect 4668 12486 4680 12538
rect 4732 12486 11372 12538
rect 11424 12486 11436 12538
rect 11488 12486 11500 12538
rect 11552 12486 11564 12538
rect 11616 12486 11628 12538
rect 11680 12486 18320 12538
rect 18372 12486 18384 12538
rect 18436 12486 18448 12538
rect 18500 12486 18512 12538
rect 18564 12486 18576 12538
rect 18628 12486 25268 12538
rect 25320 12486 25332 12538
rect 25384 12486 25396 12538
rect 25448 12486 25460 12538
rect 25512 12486 25524 12538
rect 25576 12486 28888 12538
rect 1104 12464 28888 12486
rect 15381 12427 15439 12433
rect 15381 12393 15393 12427
rect 15427 12424 15439 12427
rect 18138 12424 18144 12436
rect 15427 12396 18144 12424
rect 15427 12393 15439 12396
rect 15381 12387 15439 12393
rect 12342 12248 12348 12300
rect 12400 12288 12406 12300
rect 14185 12291 14243 12297
rect 14185 12288 14197 12291
rect 12400 12260 14197 12288
rect 12400 12248 12406 12260
rect 14185 12257 14197 12260
rect 14231 12257 14243 12291
rect 14185 12251 14243 12257
rect 5169 12223 5227 12229
rect 5169 12189 5181 12223
rect 5215 12220 5227 12223
rect 6178 12220 6184 12232
rect 5215 12192 6184 12220
rect 5215 12189 5227 12192
rect 5169 12183 5227 12189
rect 6178 12180 6184 12192
rect 6236 12180 6242 12232
rect 12526 12180 12532 12232
rect 12584 12220 12590 12232
rect 13262 12220 13268 12232
rect 12584 12192 13268 12220
rect 12584 12180 12590 12192
rect 13262 12180 13268 12192
rect 13320 12220 13326 12232
rect 14369 12223 14427 12229
rect 14369 12220 14381 12223
rect 13320 12192 14381 12220
rect 13320 12180 13326 12192
rect 14369 12189 14381 12192
rect 14415 12189 14427 12223
rect 14369 12183 14427 12189
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12220 14519 12223
rect 15396 12220 15424 12387
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 14507 12192 15424 12220
rect 14507 12189 14519 12192
rect 14461 12183 14519 12189
rect 4246 12044 4252 12096
rect 4304 12084 4310 12096
rect 4985 12087 5043 12093
rect 4985 12084 4997 12087
rect 4304 12056 4997 12084
rect 4304 12044 4310 12056
rect 4985 12053 4997 12056
rect 5031 12053 5043 12087
rect 4985 12047 5043 12053
rect 14734 12044 14740 12096
rect 14792 12084 14798 12096
rect 14829 12087 14887 12093
rect 14829 12084 14841 12087
rect 14792 12056 14841 12084
rect 14792 12044 14798 12056
rect 14829 12053 14841 12056
rect 14875 12053 14887 12087
rect 14829 12047 14887 12053
rect 1104 11994 28888 12016
rect 1104 11942 7898 11994
rect 7950 11942 7962 11994
rect 8014 11942 8026 11994
rect 8078 11942 8090 11994
rect 8142 11942 8154 11994
rect 8206 11942 14846 11994
rect 14898 11942 14910 11994
rect 14962 11942 14974 11994
rect 15026 11942 15038 11994
rect 15090 11942 15102 11994
rect 15154 11942 21794 11994
rect 21846 11942 21858 11994
rect 21910 11942 21922 11994
rect 21974 11942 21986 11994
rect 22038 11942 22050 11994
rect 22102 11942 28888 11994
rect 1104 11920 28888 11942
rect 9585 11883 9643 11889
rect 9585 11849 9597 11883
rect 9631 11880 9643 11883
rect 9858 11880 9864 11892
rect 9631 11852 9864 11880
rect 9631 11849 9643 11852
rect 9585 11843 9643 11849
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 14826 11744 14832 11756
rect 9246 11716 14832 11744
rect 14826 11704 14832 11716
rect 14884 11704 14890 11756
rect 7837 11679 7895 11685
rect 7837 11645 7849 11679
rect 7883 11645 7895 11679
rect 7837 11639 7895 11645
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11676 8171 11679
rect 11790 11676 11796 11688
rect 8159 11648 11796 11676
rect 8159 11645 8171 11648
rect 8113 11639 8171 11645
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 4617 11543 4675 11549
rect 4617 11540 4629 11543
rect 4396 11512 4629 11540
rect 4396 11500 4402 11512
rect 4617 11509 4629 11512
rect 4663 11509 4675 11543
rect 7852 11540 7880 11639
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 8478 11540 8484 11552
rect 7852 11512 8484 11540
rect 4617 11503 4675 11509
rect 8478 11500 8484 11512
rect 8536 11500 8542 11552
rect 10594 11500 10600 11552
rect 10652 11540 10658 11552
rect 10689 11543 10747 11549
rect 10689 11540 10701 11543
rect 10652 11512 10701 11540
rect 10652 11500 10658 11512
rect 10689 11509 10701 11512
rect 10735 11509 10747 11543
rect 11698 11540 11704 11552
rect 11659 11512 11704 11540
rect 10689 11503 10747 11509
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 1104 11450 28888 11472
rect 1104 11398 4424 11450
rect 4476 11398 4488 11450
rect 4540 11398 4552 11450
rect 4604 11398 4616 11450
rect 4668 11398 4680 11450
rect 4732 11398 11372 11450
rect 11424 11398 11436 11450
rect 11488 11398 11500 11450
rect 11552 11398 11564 11450
rect 11616 11398 11628 11450
rect 11680 11398 18320 11450
rect 18372 11398 18384 11450
rect 18436 11398 18448 11450
rect 18500 11398 18512 11450
rect 18564 11398 18576 11450
rect 18628 11398 25268 11450
rect 25320 11398 25332 11450
rect 25384 11398 25396 11450
rect 25448 11398 25460 11450
rect 25512 11398 25524 11450
rect 25576 11398 28888 11450
rect 1104 11376 28888 11398
rect 3142 11296 3148 11348
rect 3200 11336 3206 11348
rect 3237 11339 3295 11345
rect 3237 11336 3249 11339
rect 3200 11308 3249 11336
rect 3200 11296 3206 11308
rect 3237 11305 3249 11308
rect 3283 11305 3295 11339
rect 3237 11299 3295 11305
rect 5721 11339 5779 11345
rect 5721 11305 5733 11339
rect 5767 11336 5779 11339
rect 6362 11336 6368 11348
rect 5767 11308 6368 11336
rect 5767 11305 5779 11308
rect 5721 11299 5779 11305
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 12253 11339 12311 11345
rect 12253 11305 12265 11339
rect 12299 11336 12311 11339
rect 13630 11336 13636 11348
rect 12299 11308 13636 11336
rect 12299 11305 12311 11308
rect 12253 11299 12311 11305
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 14826 11336 14832 11348
rect 14787 11308 14832 11336
rect 14826 11296 14832 11308
rect 14884 11296 14890 11348
rect 3970 11268 3976 11280
rect 2884 11240 3976 11268
rect 1765 11203 1823 11209
rect 1765 11169 1777 11203
rect 1811 11200 1823 11203
rect 2774 11200 2780 11212
rect 1811 11172 2780 11200
rect 1811 11169 1823 11172
rect 1765 11163 1823 11169
rect 2774 11160 2780 11172
rect 2832 11160 2838 11212
rect 1486 11132 1492 11144
rect 1447 11104 1492 11132
rect 1486 11092 1492 11104
rect 1544 11092 1550 11144
rect 2884 11118 2912 11240
rect 3970 11228 3976 11240
rect 4028 11228 4034 11280
rect 4246 11200 4252 11212
rect 4207 11172 4252 11200
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 10781 11203 10839 11209
rect 10781 11169 10793 11203
rect 10827 11200 10839 11203
rect 13906 11200 13912 11212
rect 10827 11172 13912 11200
rect 10827 11169 10839 11172
rect 10781 11163 10839 11169
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 3970 11132 3976 11144
rect 3931 11104 3976 11132
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 10318 11092 10324 11144
rect 10376 11132 10382 11144
rect 10505 11135 10563 11141
rect 10505 11132 10517 11135
rect 10376 11104 10517 11132
rect 10376 11092 10382 11104
rect 10505 11101 10517 11104
rect 10551 11101 10563 11135
rect 10505 11095 10563 11101
rect 14090 11092 14096 11144
rect 14148 11132 14154 11144
rect 14642 11132 14648 11144
rect 14148 11104 14648 11132
rect 14148 11092 14154 11104
rect 14642 11092 14648 11104
rect 14700 11132 14706 11144
rect 14737 11135 14795 11141
rect 14737 11132 14749 11135
rect 14700 11104 14749 11132
rect 14700 11092 14706 11104
rect 14737 11101 14749 11104
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 4798 11024 4804 11076
rect 4856 11024 4862 11076
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 9732 11036 11270 11064
rect 9732 11024 9738 11036
rect 1104 10906 28888 10928
rect 1104 10854 7898 10906
rect 7950 10854 7962 10906
rect 8014 10854 8026 10906
rect 8078 10854 8090 10906
rect 8142 10854 8154 10906
rect 8206 10854 14846 10906
rect 14898 10854 14910 10906
rect 14962 10854 14974 10906
rect 15026 10854 15038 10906
rect 15090 10854 15102 10906
rect 15154 10854 21794 10906
rect 21846 10854 21858 10906
rect 21910 10854 21922 10906
rect 21974 10854 21986 10906
rect 22038 10854 22050 10906
rect 22102 10854 28888 10906
rect 1104 10832 28888 10854
rect 1486 10752 1492 10804
rect 1544 10792 1550 10804
rect 3970 10792 3976 10804
rect 1544 10764 3976 10792
rect 1544 10752 1550 10764
rect 1872 10665 1900 10764
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 9030 10792 9036 10804
rect 8991 10764 9036 10792
rect 9030 10752 9036 10764
rect 9088 10752 9094 10804
rect 13262 10792 13268 10804
rect 13223 10764 13268 10792
rect 13262 10752 13268 10764
rect 13320 10752 13326 10804
rect 2130 10724 2136 10736
rect 2091 10696 2136 10724
rect 2130 10684 2136 10696
rect 2188 10684 2194 10736
rect 3878 10724 3884 10736
rect 3358 10696 3884 10724
rect 3878 10684 3884 10696
rect 3936 10684 3942 10736
rect 4338 10724 4344 10736
rect 4299 10696 4344 10724
rect 4338 10684 4344 10696
rect 4396 10684 4402 10736
rect 7282 10684 7288 10736
rect 7340 10684 7346 10736
rect 9490 10684 9496 10736
rect 9548 10684 9554 10736
rect 10505 10727 10563 10733
rect 10505 10693 10517 10727
rect 10551 10724 10563 10727
rect 10778 10724 10784 10736
rect 10551 10696 10784 10724
rect 10551 10693 10563 10696
rect 10505 10687 10563 10693
rect 10778 10684 10784 10696
rect 10836 10684 10842 10736
rect 13722 10724 13728 10736
rect 13018 10696 13728 10724
rect 13722 10684 13728 10696
rect 13780 10684 13786 10736
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 5442 10616 5448 10668
rect 5500 10616 5506 10668
rect 5810 10616 5816 10668
rect 5868 10656 5874 10668
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 5868 10628 6745 10656
rect 5868 10616 5874 10628
rect 6733 10625 6745 10628
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 14734 10616 14740 10668
rect 14792 10656 14798 10668
rect 15013 10659 15071 10665
rect 15013 10656 15025 10659
rect 14792 10628 15025 10656
rect 14792 10616 14798 10628
rect 15013 10625 15025 10628
rect 15059 10625 15071 10659
rect 15013 10619 15071 10625
rect 4062 10588 4068 10600
rect 4023 10560 4068 10588
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 6362 10588 6368 10600
rect 6323 10560 6368 10588
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 6638 10548 6644 10600
rect 6696 10588 6702 10600
rect 8205 10591 8263 10597
rect 8205 10588 8217 10591
rect 6696 10560 8217 10588
rect 6696 10548 6702 10560
rect 8205 10557 8217 10560
rect 8251 10557 8263 10591
rect 10781 10591 10839 10597
rect 10781 10588 10793 10591
rect 8205 10551 8263 10557
rect 10704 10560 10793 10588
rect 3605 10455 3663 10461
rect 3605 10421 3617 10455
rect 3651 10452 3663 10455
rect 4154 10452 4160 10464
rect 3651 10424 4160 10452
rect 3651 10421 3663 10424
rect 3605 10415 3663 10421
rect 4154 10412 4160 10424
rect 4212 10412 4218 10464
rect 5810 10452 5816 10464
rect 5771 10424 5816 10452
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 10318 10412 10324 10464
rect 10376 10452 10382 10464
rect 10704 10452 10732 10560
rect 10781 10557 10793 10560
rect 10827 10588 10839 10591
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 10827 10560 11529 10588
rect 10827 10557 10839 10560
rect 10781 10551 10839 10557
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 11793 10591 11851 10597
rect 11793 10557 11805 10591
rect 11839 10588 11851 10591
rect 11839 10560 14872 10588
rect 11839 10557 11851 10560
rect 11793 10551 11851 10557
rect 14844 10529 14872 10560
rect 14829 10523 14887 10529
rect 14829 10489 14841 10523
rect 14875 10489 14887 10523
rect 14829 10483 14887 10489
rect 10376 10424 10732 10452
rect 10376 10412 10382 10424
rect 1104 10362 28888 10384
rect 1104 10310 4424 10362
rect 4476 10310 4488 10362
rect 4540 10310 4552 10362
rect 4604 10310 4616 10362
rect 4668 10310 4680 10362
rect 4732 10310 11372 10362
rect 11424 10310 11436 10362
rect 11488 10310 11500 10362
rect 11552 10310 11564 10362
rect 11616 10310 11628 10362
rect 11680 10310 18320 10362
rect 18372 10310 18384 10362
rect 18436 10310 18448 10362
rect 18500 10310 18512 10362
rect 18564 10310 18576 10362
rect 18628 10310 25268 10362
rect 25320 10310 25332 10362
rect 25384 10310 25396 10362
rect 25448 10310 25460 10362
rect 25512 10310 25524 10362
rect 25576 10310 28888 10362
rect 1104 10288 28888 10310
rect 3234 10248 3240 10260
rect 3195 10220 3240 10248
rect 3234 10208 3240 10220
rect 3292 10208 3298 10260
rect 5810 10208 5816 10260
rect 5868 10248 5874 10260
rect 13998 10248 14004 10260
rect 5868 10220 14004 10248
rect 5868 10208 5874 10220
rect 13998 10208 14004 10220
rect 14056 10208 14062 10260
rect 7374 10140 7380 10192
rect 7432 10180 7438 10192
rect 7975 10183 8033 10189
rect 7975 10180 7987 10183
rect 7432 10152 7987 10180
rect 7432 10140 7438 10152
rect 7975 10149 7987 10152
rect 8021 10149 8033 10183
rect 7975 10143 8033 10149
rect 1762 10112 1768 10124
rect 1723 10084 1768 10112
rect 1762 10072 1768 10084
rect 1820 10072 1826 10124
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10112 6239 10115
rect 6362 10112 6368 10124
rect 6227 10084 6368 10112
rect 6227 10081 6239 10084
rect 6181 10075 6239 10081
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 6549 10115 6607 10121
rect 6549 10112 6561 10115
rect 6512 10084 6561 10112
rect 6512 10072 6518 10084
rect 6549 10081 6561 10084
rect 6595 10081 6607 10115
rect 10594 10112 10600 10124
rect 10555 10084 10600 10112
rect 6549 10075 6607 10081
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 11146 10072 11152 10124
rect 11204 10112 11210 10124
rect 14553 10115 14611 10121
rect 14553 10112 14565 10115
rect 11204 10084 14565 10112
rect 11204 10072 11210 10084
rect 14553 10081 14565 10084
rect 14599 10081 14611 10115
rect 14553 10075 14611 10081
rect 1486 10044 1492 10056
rect 1447 10016 1492 10044
rect 1486 10004 1492 10016
rect 1544 10004 1550 10056
rect 10318 10044 10324 10056
rect 10279 10016 10324 10044
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 14642 10044 14648 10056
rect 14603 10016 14648 10044
rect 14642 10004 14648 10016
rect 14700 10004 14706 10056
rect 3510 9976 3516 9988
rect 2990 9948 3516 9976
rect 3510 9936 3516 9948
rect 3568 9936 3574 9988
rect 6914 9936 6920 9988
rect 6972 9936 6978 9988
rect 12710 9976 12716 9988
rect 11822 9948 12716 9976
rect 12710 9936 12716 9948
rect 12768 9936 12774 9988
rect 12069 9911 12127 9917
rect 12069 9877 12081 9911
rect 12115 9908 12127 9911
rect 13722 9908 13728 9920
rect 12115 9880 13728 9908
rect 12115 9877 12127 9880
rect 12069 9871 12127 9877
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 1104 9818 28888 9840
rect 1104 9766 7898 9818
rect 7950 9766 7962 9818
rect 8014 9766 8026 9818
rect 8078 9766 8090 9818
rect 8142 9766 8154 9818
rect 8206 9766 14846 9818
rect 14898 9766 14910 9818
rect 14962 9766 14974 9818
rect 15026 9766 15038 9818
rect 15090 9766 15102 9818
rect 15154 9766 21794 9818
rect 21846 9766 21858 9818
rect 21910 9766 21922 9818
rect 21974 9766 21986 9818
rect 22038 9766 22050 9818
rect 22102 9766 28888 9818
rect 1104 9744 28888 9766
rect 2038 9636 2044 9648
rect 1999 9608 2044 9636
rect 2038 9596 2044 9608
rect 2096 9596 2102 9648
rect 4982 9636 4988 9648
rect 3266 9608 4988 9636
rect 4982 9596 4988 9608
rect 5040 9596 5046 9648
rect 11146 9636 11152 9648
rect 7682 9608 11152 9636
rect 11146 9596 11152 9608
rect 11204 9596 11210 9648
rect 11698 9596 11704 9648
rect 11756 9636 11762 9648
rect 11793 9639 11851 9645
rect 11793 9636 11805 9639
rect 11756 9608 11805 9636
rect 11756 9596 11762 9608
rect 11793 9605 11805 9608
rect 11839 9605 11851 9639
rect 11793 9599 11851 9605
rect 13722 9596 13728 9648
rect 13780 9636 13786 9648
rect 13780 9608 14136 9636
rect 13780 9596 13786 9608
rect 8389 9571 8447 9577
rect 8389 9537 8401 9571
rect 8435 9568 8447 9571
rect 8478 9568 8484 9580
rect 8435 9540 8484 9568
rect 8435 9537 8447 9540
rect 8389 9531 8447 9537
rect 8478 9528 8484 9540
rect 8536 9568 8542 9580
rect 10318 9568 10324 9580
rect 8536 9540 10324 9568
rect 8536 9528 8542 9540
rect 10318 9528 10324 9540
rect 10376 9568 10382 9580
rect 14108 9577 14136 9608
rect 14642 9596 14648 9648
rect 14700 9636 14706 9648
rect 14700 9608 16574 9636
rect 14700 9596 14706 9608
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 10376 9540 11529 9568
rect 10376 9528 10382 9540
rect 11517 9537 11529 9540
rect 11563 9537 11575 9571
rect 14001 9571 14059 9577
rect 11517 9531 11575 9537
rect 1486 9460 1492 9512
rect 1544 9500 1550 9512
rect 1765 9503 1823 9509
rect 1765 9500 1777 9503
rect 1544 9472 1777 9500
rect 1544 9460 1550 9472
rect 1765 9469 1777 9472
rect 1811 9469 1823 9503
rect 1765 9463 1823 9469
rect 1780 9364 1808 9463
rect 3326 9460 3332 9512
rect 3384 9500 3390 9512
rect 3513 9503 3571 9509
rect 3513 9500 3525 9503
rect 3384 9472 3525 9500
rect 3384 9460 3390 9472
rect 3513 9469 3525 9472
rect 3559 9469 3571 9503
rect 3513 9463 3571 9469
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 6641 9503 6699 9509
rect 6641 9500 6653 9503
rect 6604 9472 6653 9500
rect 6604 9460 6610 9472
rect 6641 9469 6653 9472
rect 6687 9469 6699 9503
rect 6641 9463 6699 9469
rect 7742 9460 7748 9512
rect 7800 9500 7806 9512
rect 8113 9503 8171 9509
rect 8113 9500 8125 9503
rect 7800 9472 8125 9500
rect 7800 9460 7806 9472
rect 8113 9469 8125 9472
rect 8159 9469 8171 9503
rect 8113 9463 8171 9469
rect 10686 9460 10692 9512
rect 10744 9500 10750 9512
rect 12912 9500 12940 9554
rect 14001 9537 14013 9571
rect 14047 9537 14059 9571
rect 14001 9531 14059 9537
rect 14093 9571 14151 9577
rect 14093 9537 14105 9571
rect 14139 9537 14151 9571
rect 15286 9568 15292 9580
rect 15247 9540 15292 9568
rect 14093 9531 14151 9537
rect 10744 9472 12940 9500
rect 13265 9503 13323 9509
rect 10744 9460 10750 9472
rect 13265 9469 13277 9503
rect 13311 9500 13323 9503
rect 14016 9500 14044 9531
rect 15286 9528 15292 9540
rect 15344 9528 15350 9580
rect 16546 9568 16574 9608
rect 19061 9571 19119 9577
rect 19061 9568 19073 9571
rect 16546 9540 19073 9568
rect 19061 9537 19073 9540
rect 19107 9568 19119 9571
rect 19521 9571 19579 9577
rect 19521 9568 19533 9571
rect 19107 9540 19533 9568
rect 19107 9537 19119 9540
rect 19061 9531 19119 9537
rect 19521 9537 19533 9540
rect 19567 9537 19579 9571
rect 19521 9531 19579 9537
rect 13311 9472 14044 9500
rect 13311 9469 13323 9472
rect 13265 9463 13323 9469
rect 14274 9460 14280 9512
rect 14332 9500 14338 9512
rect 15013 9503 15071 9509
rect 15013 9500 15025 9503
rect 14332 9472 15025 9500
rect 14332 9460 14338 9472
rect 15013 9469 15025 9472
rect 15059 9500 15071 9503
rect 15059 9472 15516 9500
rect 15059 9469 15071 9472
rect 15013 9463 15071 9469
rect 3234 9364 3240 9376
rect 1780 9336 3240 9364
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 13998 9364 14004 9376
rect 13959 9336 14004 9364
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 14369 9367 14427 9373
rect 14369 9333 14381 9367
rect 14415 9364 14427 9367
rect 15378 9364 15384 9376
rect 14415 9336 15384 9364
rect 14415 9333 14427 9336
rect 14369 9327 14427 9333
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 15488 9364 15516 9472
rect 16666 9364 16672 9376
rect 15488 9336 16672 9364
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 18966 9364 18972 9376
rect 18927 9336 18972 9364
rect 18966 9324 18972 9336
rect 19024 9324 19030 9376
rect 19610 9364 19616 9376
rect 19571 9336 19616 9364
rect 19610 9324 19616 9336
rect 19668 9324 19674 9376
rect 1104 9274 28888 9296
rect 1104 9222 4424 9274
rect 4476 9222 4488 9274
rect 4540 9222 4552 9274
rect 4604 9222 4616 9274
rect 4668 9222 4680 9274
rect 4732 9222 11372 9274
rect 11424 9222 11436 9274
rect 11488 9222 11500 9274
rect 11552 9222 11564 9274
rect 11616 9222 11628 9274
rect 11680 9222 18320 9274
rect 18372 9222 18384 9274
rect 18436 9222 18448 9274
rect 18500 9222 18512 9274
rect 18564 9222 18576 9274
rect 18628 9222 25268 9274
rect 25320 9222 25332 9274
rect 25384 9222 25396 9274
rect 25448 9222 25460 9274
rect 25512 9222 25524 9274
rect 25576 9222 28888 9274
rect 1104 9200 28888 9222
rect 7558 9120 7564 9172
rect 7616 9160 7622 9172
rect 7745 9163 7803 9169
rect 7745 9160 7757 9163
rect 7616 9132 7757 9160
rect 7616 9120 7622 9132
rect 7745 9129 7757 9132
rect 7791 9129 7803 9163
rect 7745 9123 7803 9129
rect 12710 9120 12716 9172
rect 12768 9160 12774 9172
rect 14369 9163 14427 9169
rect 14369 9160 14381 9163
rect 12768 9132 14381 9160
rect 12768 9120 12774 9132
rect 14369 9129 14381 9132
rect 14415 9129 14427 9163
rect 19610 9160 19616 9172
rect 14369 9123 14427 9129
rect 16546 9132 19616 9160
rect 3234 8984 3240 9036
rect 3292 9024 3298 9036
rect 4062 9024 4068 9036
rect 3292 8996 4068 9024
rect 3292 8984 3298 8996
rect 4062 8984 4068 8996
rect 4120 9024 4126 9036
rect 5997 9027 6055 9033
rect 5997 9024 6009 9027
rect 4120 8996 6009 9024
rect 4120 8984 4126 8996
rect 5997 8993 6009 8996
rect 6043 9024 6055 9027
rect 6362 9024 6368 9036
rect 6043 8996 6368 9024
rect 6043 8993 6055 8996
rect 5997 8987 6055 8993
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 6638 8984 6644 9036
rect 6696 9024 6702 9036
rect 7006 9024 7012 9036
rect 6696 8996 7012 9024
rect 6696 8984 6702 8996
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 7558 8984 7564 9036
rect 7616 9024 7622 9036
rect 16546 9024 16574 9132
rect 19610 9120 19616 9132
rect 19668 9120 19674 9172
rect 7616 8996 16574 9024
rect 7616 8984 7622 8996
rect 10042 8956 10048 8968
rect 10003 8928 10048 8956
rect 10042 8916 10048 8928
rect 10100 8916 10106 8968
rect 14461 8959 14519 8965
rect 14461 8925 14473 8959
rect 14507 8956 14519 8959
rect 14734 8956 14740 8968
rect 14507 8928 14740 8956
rect 14507 8925 14519 8928
rect 14461 8919 14519 8925
rect 14734 8916 14740 8928
rect 14792 8916 14798 8968
rect 6273 8891 6331 8897
rect 6273 8857 6285 8891
rect 6319 8888 6331 8891
rect 6546 8888 6552 8900
rect 6319 8860 6552 8888
rect 6319 8857 6331 8860
rect 6273 8851 6331 8857
rect 6546 8848 6552 8860
rect 6604 8848 6610 8900
rect 7650 8888 7656 8900
rect 7498 8860 7656 8888
rect 7650 8848 7656 8860
rect 7708 8848 7714 8900
rect 1104 8730 28888 8752
rect 1104 8678 7898 8730
rect 7950 8678 7962 8730
rect 8014 8678 8026 8730
rect 8078 8678 8090 8730
rect 8142 8678 8154 8730
rect 8206 8678 14846 8730
rect 14898 8678 14910 8730
rect 14962 8678 14974 8730
rect 15026 8678 15038 8730
rect 15090 8678 15102 8730
rect 15154 8678 21794 8730
rect 21846 8678 21858 8730
rect 21910 8678 21922 8730
rect 21974 8678 21986 8730
rect 22038 8678 22050 8730
rect 22102 8678 28888 8730
rect 1104 8656 28888 8678
rect 4798 8548 4804 8560
rect 4738 8520 4804 8548
rect 4798 8508 4804 8520
rect 4856 8508 4862 8560
rect 9493 8551 9551 8557
rect 9493 8517 9505 8551
rect 9539 8548 9551 8551
rect 9766 8548 9772 8560
rect 9539 8520 9772 8548
rect 9539 8517 9551 8520
rect 9493 8511 9551 8517
rect 9766 8508 9772 8520
rect 9824 8508 9830 8560
rect 12342 8548 12348 8560
rect 10718 8520 12348 8548
rect 12342 8508 12348 8520
rect 12400 8508 12406 8560
rect 3234 8480 3240 8492
rect 3195 8452 3240 8480
rect 3234 8440 3240 8452
rect 3292 8440 3298 8492
rect 8478 8440 8484 8492
rect 8536 8480 8542 8492
rect 9217 8483 9275 8489
rect 9217 8480 9229 8483
rect 8536 8452 9229 8480
rect 8536 8440 8542 8452
rect 9217 8449 9229 8452
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8480 14151 8483
rect 14734 8480 14740 8492
rect 14139 8452 14740 8480
rect 14139 8449 14151 8452
rect 14093 8443 14151 8449
rect 14734 8440 14740 8452
rect 14792 8440 14798 8492
rect 3510 8412 3516 8424
rect 3471 8384 3516 8412
rect 3510 8372 3516 8384
rect 3568 8372 3574 8424
rect 13998 8412 14004 8424
rect 13959 8384 14004 8412
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 4985 8347 5043 8353
rect 4985 8313 4997 8347
rect 5031 8344 5043 8347
rect 6270 8344 6276 8356
rect 5031 8316 6276 8344
rect 5031 8313 5043 8316
rect 4985 8307 5043 8313
rect 6270 8304 6276 8316
rect 6328 8304 6334 8356
rect 6638 8304 6644 8356
rect 6696 8344 6702 8356
rect 7101 8347 7159 8353
rect 7101 8344 7113 8347
rect 6696 8316 7113 8344
rect 6696 8304 6702 8316
rect 7101 8313 7113 8316
rect 7147 8313 7159 8347
rect 7101 8307 7159 8313
rect 10965 8347 11023 8353
rect 10965 8313 10977 8347
rect 11011 8344 11023 8347
rect 14090 8344 14096 8356
rect 11011 8316 14096 8344
rect 11011 8313 11023 8316
rect 10965 8307 11023 8313
rect 14090 8304 14096 8316
rect 14148 8304 14154 8356
rect 11238 8236 11244 8288
rect 11296 8276 11302 8288
rect 11517 8279 11575 8285
rect 11517 8276 11529 8279
rect 11296 8248 11529 8276
rect 11296 8236 11302 8248
rect 11517 8245 11529 8248
rect 11563 8245 11575 8279
rect 11517 8239 11575 8245
rect 1104 8186 28888 8208
rect 1104 8134 4424 8186
rect 4476 8134 4488 8186
rect 4540 8134 4552 8186
rect 4604 8134 4616 8186
rect 4668 8134 4680 8186
rect 4732 8134 11372 8186
rect 11424 8134 11436 8186
rect 11488 8134 11500 8186
rect 11552 8134 11564 8186
rect 11616 8134 11628 8186
rect 11680 8134 18320 8186
rect 18372 8134 18384 8186
rect 18436 8134 18448 8186
rect 18500 8134 18512 8186
rect 18564 8134 18576 8186
rect 18628 8134 25268 8186
rect 25320 8134 25332 8186
rect 25384 8134 25396 8186
rect 25448 8134 25460 8186
rect 25512 8134 25524 8186
rect 25576 8134 28888 8186
rect 1104 8112 28888 8134
rect 3510 8032 3516 8084
rect 3568 8072 3574 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 3568 8044 3801 8072
rect 3568 8032 3574 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 9766 8072 9772 8084
rect 9727 8044 9772 8072
rect 3789 8035 3847 8041
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 12342 8032 12348 8084
rect 12400 8072 12406 8084
rect 13449 8075 13507 8081
rect 13449 8072 13461 8075
rect 12400 8044 13461 8072
rect 12400 8032 12406 8044
rect 13449 8041 13461 8044
rect 13495 8041 13507 8075
rect 14090 8072 14096 8084
rect 14051 8044 14096 8072
rect 13449 8035 13507 8041
rect 14090 8032 14096 8044
rect 14148 8032 14154 8084
rect 14553 8075 14611 8081
rect 14553 8041 14565 8075
rect 14599 8072 14611 8075
rect 15197 8075 15255 8081
rect 15197 8072 15209 8075
rect 14599 8044 15209 8072
rect 14599 8041 14611 8044
rect 14553 8035 14611 8041
rect 15197 8041 15209 8044
rect 15243 8041 15255 8075
rect 15562 8072 15568 8084
rect 15523 8044 15568 8072
rect 15197 8035 15255 8041
rect 15562 8032 15568 8044
rect 15620 8032 15626 8084
rect 1489 7939 1547 7945
rect 1489 7905 1501 7939
rect 1535 7936 1547 7939
rect 3234 7936 3240 7948
rect 1535 7908 3240 7936
rect 1535 7905 1547 7908
rect 1489 7899 1547 7905
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 8389 7939 8447 7945
rect 8389 7905 8401 7939
rect 8435 7936 8447 7939
rect 8478 7936 8484 7948
rect 8435 7908 8484 7936
rect 8435 7905 8447 7908
rect 8389 7899 8447 7905
rect 8478 7896 8484 7908
rect 8536 7936 8542 7948
rect 10597 7939 10655 7945
rect 10597 7936 10609 7939
rect 8536 7908 10609 7936
rect 8536 7896 8542 7908
rect 10597 7905 10609 7908
rect 10643 7905 10655 7939
rect 10597 7899 10655 7905
rect 10873 7939 10931 7945
rect 10873 7905 10885 7939
rect 10919 7936 10931 7939
rect 11238 7936 11244 7948
rect 10919 7908 11244 7936
rect 10919 7905 10931 7908
rect 10873 7899 10931 7905
rect 11238 7896 11244 7908
rect 11296 7896 11302 7948
rect 11330 7896 11336 7948
rect 11388 7936 11394 7948
rect 14185 7939 14243 7945
rect 14185 7936 14197 7939
rect 11388 7908 14197 7936
rect 11388 7896 11394 7908
rect 14185 7905 14197 7908
rect 14231 7905 14243 7939
rect 14185 7899 14243 7905
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7868 13599 7871
rect 13587 7840 14228 7868
rect 13587 7837 13599 7840
rect 13541 7831 13599 7837
rect 1762 7800 1768 7812
rect 1723 7772 1768 7800
rect 1762 7760 1768 7772
rect 1820 7760 1826 7812
rect 3694 7800 3700 7812
rect 2990 7772 3700 7800
rect 3694 7760 3700 7772
rect 3752 7760 3758 7812
rect 4338 7760 4344 7812
rect 4396 7800 4402 7812
rect 6641 7803 6699 7809
rect 6641 7800 6653 7803
rect 4396 7772 6653 7800
rect 4396 7760 4402 7772
rect 6641 7769 6653 7772
rect 6687 7800 6699 7803
rect 7650 7800 7656 7812
rect 6687 7772 7656 7800
rect 6687 7769 6699 7772
rect 6641 7763 6699 7769
rect 7650 7760 7656 7772
rect 7708 7760 7714 7812
rect 12250 7800 12256 7812
rect 12098 7772 12256 7800
rect 12250 7760 12256 7772
rect 12308 7760 12314 7812
rect 14093 7803 14151 7809
rect 14093 7800 14105 7803
rect 12360 7772 14105 7800
rect 3237 7735 3295 7741
rect 3237 7701 3249 7735
rect 3283 7732 3295 7735
rect 4890 7732 4896 7744
rect 3283 7704 4896 7732
rect 3283 7701 3295 7704
rect 3237 7695 3295 7701
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 6178 7732 6184 7744
rect 6139 7704 6184 7732
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 12360 7741 12388 7772
rect 14093 7769 14105 7772
rect 14139 7769 14151 7803
rect 14200 7800 14228 7840
rect 14274 7828 14280 7880
rect 14332 7868 14338 7880
rect 14369 7871 14427 7877
rect 14369 7868 14381 7871
rect 14332 7840 14381 7868
rect 14332 7828 14338 7840
rect 14369 7837 14381 7840
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 14458 7828 14464 7880
rect 14516 7868 14522 7880
rect 15197 7871 15255 7877
rect 15197 7868 15209 7871
rect 14516 7840 15209 7868
rect 14516 7828 14522 7840
rect 15197 7837 15209 7840
rect 15243 7837 15255 7871
rect 15378 7868 15384 7880
rect 15339 7840 15384 7868
rect 15197 7831 15255 7837
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 14734 7800 14740 7812
rect 14200 7772 14740 7800
rect 14093 7763 14151 7769
rect 14734 7760 14740 7772
rect 14792 7800 14798 7812
rect 16485 7803 16543 7809
rect 16485 7800 16497 7803
rect 14792 7772 16497 7800
rect 14792 7760 14798 7772
rect 16485 7769 16497 7772
rect 16531 7769 16543 7803
rect 16485 7763 16543 7769
rect 16666 7760 16672 7812
rect 16724 7800 16730 7812
rect 16724 7772 16817 7800
rect 16724 7760 16730 7772
rect 12345 7735 12403 7741
rect 12345 7701 12357 7735
rect 12391 7701 12403 7735
rect 16684 7732 16712 7760
rect 17313 7735 17371 7741
rect 17313 7732 17325 7735
rect 16684 7704 17325 7732
rect 12345 7695 12403 7701
rect 17313 7701 17325 7704
rect 17359 7732 17371 7735
rect 23290 7732 23296 7744
rect 17359 7704 23296 7732
rect 17359 7701 17371 7704
rect 17313 7695 17371 7701
rect 23290 7692 23296 7704
rect 23348 7692 23354 7744
rect 1104 7642 28888 7664
rect 1104 7590 7898 7642
rect 7950 7590 7962 7642
rect 8014 7590 8026 7642
rect 8078 7590 8090 7642
rect 8142 7590 8154 7642
rect 8206 7590 14846 7642
rect 14898 7590 14910 7642
rect 14962 7590 14974 7642
rect 15026 7590 15038 7642
rect 15090 7590 15102 7642
rect 15154 7590 21794 7642
rect 21846 7590 21858 7642
rect 21910 7590 21922 7642
rect 21974 7590 21986 7642
rect 22038 7590 22050 7642
rect 22102 7590 28888 7642
rect 1104 7568 28888 7590
rect 3053 7531 3111 7537
rect 3053 7497 3065 7531
rect 3099 7528 3111 7531
rect 3234 7528 3240 7540
rect 3099 7500 3240 7528
rect 3099 7497 3111 7500
rect 3053 7491 3111 7497
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 10965 7531 11023 7537
rect 10965 7497 10977 7531
rect 11011 7528 11023 7531
rect 11330 7528 11336 7540
rect 11011 7500 11336 7528
rect 11011 7497 11023 7500
rect 10965 7491 11023 7497
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 12250 7488 12256 7540
rect 12308 7528 12314 7540
rect 14093 7531 14151 7537
rect 14093 7528 14105 7531
rect 12308 7500 14105 7528
rect 12308 7488 12314 7500
rect 14093 7497 14105 7500
rect 14139 7497 14151 7531
rect 14093 7491 14151 7497
rect 6178 7420 6184 7472
rect 6236 7460 6242 7472
rect 6733 7463 6791 7469
rect 6733 7460 6745 7463
rect 6236 7432 6745 7460
rect 6236 7420 6242 7432
rect 6733 7429 6745 7432
rect 6779 7429 6791 7463
rect 13998 7460 14004 7472
rect 10718 7432 14004 7460
rect 6733 7423 6791 7429
rect 13998 7420 14004 7432
rect 14056 7420 14062 7472
rect 1762 7352 1768 7404
rect 1820 7392 1826 7404
rect 1949 7395 2007 7401
rect 1949 7392 1961 7395
rect 1820 7364 1961 7392
rect 1820 7352 1826 7364
rect 1949 7361 1961 7364
rect 1995 7361 2007 7395
rect 4338 7392 4344 7404
rect 4299 7364 4344 7392
rect 1949 7355 2007 7361
rect 4338 7352 4344 7364
rect 4396 7352 4402 7404
rect 8478 7352 8484 7404
rect 8536 7392 8542 7404
rect 9217 7395 9275 7401
rect 9217 7392 9229 7395
rect 8536 7364 9229 7392
rect 8536 7352 8542 7364
rect 9217 7361 9229 7364
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 13541 7395 13599 7401
rect 13541 7361 13553 7395
rect 13587 7361 13599 7395
rect 13541 7355 13599 7361
rect 14185 7395 14243 7401
rect 14185 7361 14197 7395
rect 14231 7392 14243 7395
rect 14734 7392 14740 7404
rect 14231 7364 14740 7392
rect 14231 7361 14243 7364
rect 14185 7355 14243 7361
rect 9493 7327 9551 7333
rect 9493 7293 9505 7327
rect 9539 7324 9551 7327
rect 10042 7324 10048 7336
rect 9539 7296 10048 7324
rect 9539 7293 9551 7296
rect 9493 7287 9551 7293
rect 10042 7284 10048 7296
rect 10100 7284 10106 7336
rect 13556 7324 13584 7355
rect 14734 7352 14740 7364
rect 14792 7392 14798 7404
rect 14829 7395 14887 7401
rect 14829 7392 14841 7395
rect 14792 7364 14841 7392
rect 14792 7352 14798 7364
rect 14829 7361 14841 7364
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 14642 7324 14648 7336
rect 13556 7296 14648 7324
rect 14642 7284 14648 7296
rect 14700 7284 14706 7336
rect 10778 7216 10784 7268
rect 10836 7256 10842 7268
rect 13449 7259 13507 7265
rect 13449 7256 13461 7259
rect 10836 7228 13461 7256
rect 10836 7216 10842 7228
rect 13449 7225 13461 7228
rect 13495 7225 13507 7259
rect 13449 7219 13507 7225
rect 4982 7188 4988 7200
rect 4943 7160 4988 7188
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 5810 7188 5816 7200
rect 5771 7160 5816 7188
rect 5810 7148 5816 7160
rect 5868 7148 5874 7200
rect 7650 7148 7656 7200
rect 7708 7188 7714 7200
rect 8021 7191 8079 7197
rect 8021 7188 8033 7191
rect 7708 7160 8033 7188
rect 7708 7148 7714 7160
rect 8021 7157 8033 7160
rect 8067 7157 8079 7191
rect 8021 7151 8079 7157
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 14737 7191 14795 7197
rect 14737 7188 14749 7191
rect 13228 7160 14749 7188
rect 13228 7148 13234 7160
rect 14737 7157 14749 7160
rect 14783 7157 14795 7191
rect 14737 7151 14795 7157
rect 1104 7098 28888 7120
rect 1104 7046 4424 7098
rect 4476 7046 4488 7098
rect 4540 7046 4552 7098
rect 4604 7046 4616 7098
rect 4668 7046 4680 7098
rect 4732 7046 11372 7098
rect 11424 7046 11436 7098
rect 11488 7046 11500 7098
rect 11552 7046 11564 7098
rect 11616 7046 11628 7098
rect 11680 7046 18320 7098
rect 18372 7046 18384 7098
rect 18436 7046 18448 7098
rect 18500 7046 18512 7098
rect 18564 7046 18576 7098
rect 18628 7046 25268 7098
rect 25320 7046 25332 7098
rect 25384 7046 25396 7098
rect 25448 7046 25460 7098
rect 25512 7046 25524 7098
rect 25576 7046 28888 7098
rect 1104 7024 28888 7046
rect 4420 6987 4478 6993
rect 4420 6953 4432 6987
rect 4466 6984 4478 6987
rect 4982 6984 4988 6996
rect 4466 6956 4988 6984
rect 4466 6953 4478 6956
rect 4420 6947 4478 6953
rect 4982 6944 4988 6956
rect 5040 6944 5046 6996
rect 5810 6944 5816 6996
rect 5868 6984 5874 6996
rect 6622 6987 6680 6993
rect 6622 6984 6634 6987
rect 5868 6956 6634 6984
rect 5868 6944 5874 6956
rect 6622 6953 6634 6956
rect 6668 6953 6680 6987
rect 14090 6984 14096 6996
rect 14051 6956 14096 6984
rect 6622 6947 6680 6953
rect 14090 6944 14096 6956
rect 14148 6944 14154 6996
rect 4157 6851 4215 6857
rect 4157 6817 4169 6851
rect 4203 6848 4215 6851
rect 4203 6820 6408 6848
rect 4203 6817 4215 6820
rect 4157 6811 4215 6817
rect 6380 6792 6408 6820
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 10778 6848 10784 6860
rect 6788 6820 10784 6848
rect 6788 6808 6794 6820
rect 10778 6808 10784 6820
rect 10836 6808 10842 6860
rect 11238 6808 11244 6860
rect 11296 6848 11302 6860
rect 14185 6851 14243 6857
rect 14185 6848 14197 6851
rect 11296 6820 14197 6848
rect 11296 6808 11302 6820
rect 14185 6817 14197 6820
rect 14231 6817 14243 6851
rect 14185 6811 14243 6817
rect 2314 6780 2320 6792
rect 2275 6752 2320 6780
rect 2314 6740 2320 6752
rect 2372 6740 2378 6792
rect 3142 6780 3148 6792
rect 3055 6752 3148 6780
rect 3142 6740 3148 6752
rect 3200 6780 3206 6792
rect 3602 6780 3608 6792
rect 3200 6752 3608 6780
rect 3200 6740 3206 6752
rect 3602 6740 3608 6752
rect 3660 6740 3666 6792
rect 6362 6780 6368 6792
rect 6323 6752 6368 6780
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 10318 6740 10324 6792
rect 10376 6780 10382 6792
rect 10873 6783 10931 6789
rect 10873 6780 10885 6783
rect 10376 6752 10885 6780
rect 10376 6740 10382 6752
rect 10873 6749 10885 6752
rect 10919 6749 10931 6783
rect 14366 6780 14372 6792
rect 14327 6752 14372 6780
rect 10873 6743 10931 6749
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 15194 6740 15200 6792
rect 15252 6780 15258 6792
rect 16485 6783 16543 6789
rect 16485 6780 16497 6783
rect 15252 6752 16497 6780
rect 15252 6740 15258 6752
rect 16485 6749 16497 6752
rect 16531 6749 16543 6783
rect 16485 6743 16543 6749
rect 1857 6715 1915 6721
rect 1857 6681 1869 6715
rect 1903 6712 1915 6715
rect 3160 6712 3188 6740
rect 6730 6712 6736 6724
rect 1903 6684 3188 6712
rect 5658 6684 6736 6712
rect 1903 6681 1915 6684
rect 1857 6675 1915 6681
rect 6730 6672 6736 6684
rect 6788 6672 6794 6724
rect 10686 6712 10692 6724
rect 7866 6684 10692 6712
rect 10686 6672 10692 6684
rect 10744 6672 10750 6724
rect 11146 6712 11152 6724
rect 11107 6684 11152 6712
rect 11146 6672 11152 6684
rect 11204 6672 11210 6724
rect 13170 6712 13176 6724
rect 12374 6684 13176 6712
rect 13170 6672 13176 6684
rect 13228 6672 13234 6724
rect 14090 6712 14096 6724
rect 14051 6684 14096 6712
rect 14090 6672 14096 6684
rect 14148 6672 14154 6724
rect 3050 6644 3056 6656
rect 3011 6616 3056 6644
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 5902 6644 5908 6656
rect 5863 6616 5908 6644
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 6546 6604 6552 6656
rect 6604 6644 6610 6656
rect 8113 6647 8171 6653
rect 8113 6644 8125 6647
rect 6604 6616 8125 6644
rect 6604 6604 6610 6616
rect 8113 6613 8125 6616
rect 8159 6613 8171 6647
rect 8113 6607 8171 6613
rect 12621 6647 12679 6653
rect 12621 6613 12633 6647
rect 12667 6644 12679 6647
rect 12802 6644 12808 6656
rect 12667 6616 12808 6644
rect 12667 6613 12679 6616
rect 12621 6607 12679 6613
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 14550 6644 14556 6656
rect 14511 6616 14556 6644
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 16574 6604 16580 6656
rect 16632 6644 16638 6656
rect 16632 6616 16677 6644
rect 16632 6604 16638 6616
rect 1104 6554 28888 6576
rect 1104 6502 7898 6554
rect 7950 6502 7962 6554
rect 8014 6502 8026 6554
rect 8078 6502 8090 6554
rect 8142 6502 8154 6554
rect 8206 6502 14846 6554
rect 14898 6502 14910 6554
rect 14962 6502 14974 6554
rect 15026 6502 15038 6554
rect 15090 6502 15102 6554
rect 15154 6502 21794 6554
rect 21846 6502 21858 6554
rect 21910 6502 21922 6554
rect 21974 6502 21986 6554
rect 22038 6502 22050 6554
rect 22102 6502 28888 6554
rect 1104 6480 28888 6502
rect 4709 6443 4767 6449
rect 4709 6409 4721 6443
rect 4755 6440 4767 6443
rect 4798 6440 4804 6452
rect 4755 6412 4804 6440
rect 4755 6409 4767 6412
rect 4709 6403 4767 6409
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 8113 6443 8171 6449
rect 8113 6409 8125 6443
rect 8159 6440 8171 6443
rect 11238 6440 11244 6452
rect 8159 6412 11244 6440
rect 8159 6409 8171 6412
rect 8113 6403 8171 6409
rect 11238 6400 11244 6412
rect 11296 6400 11302 6452
rect 13265 6443 13323 6449
rect 13265 6409 13277 6443
rect 13311 6409 13323 6443
rect 14182 6440 14188 6452
rect 14143 6412 14188 6440
rect 13265 6403 13323 6409
rect 2314 6372 2320 6384
rect 2275 6344 2320 6372
rect 2314 6332 2320 6344
rect 2372 6332 2378 6384
rect 3602 6332 3608 6384
rect 3660 6372 3666 6384
rect 5350 6372 5356 6384
rect 3660 6344 5356 6372
rect 3660 6332 3666 6344
rect 3418 6264 3424 6316
rect 3476 6264 3482 6316
rect 4816 6313 4844 6344
rect 5350 6332 5356 6344
rect 5408 6332 5414 6384
rect 6638 6372 6644 6384
rect 6599 6344 6644 6372
rect 6638 6332 6644 6344
rect 6696 6332 6702 6384
rect 12802 6372 12808 6384
rect 12763 6344 12808 6372
rect 12802 6332 12808 6344
rect 12860 6332 12866 6384
rect 13280 6372 13308 6403
rect 14182 6400 14188 6412
rect 14240 6400 14246 6452
rect 14642 6400 14648 6452
rect 14700 6440 14706 6452
rect 14829 6443 14887 6449
rect 14829 6440 14841 6443
rect 14700 6412 14841 6440
rect 14700 6400 14706 6412
rect 14829 6409 14841 6412
rect 14875 6409 14887 6443
rect 14829 6403 14887 6409
rect 14458 6372 14464 6384
rect 13280 6344 14464 6372
rect 14458 6332 14464 6344
rect 14516 6332 14522 6384
rect 4801 6307 4859 6313
rect 4801 6273 4813 6307
rect 4847 6273 4859 6307
rect 4801 6267 4859 6273
rect 7742 6264 7748 6316
rect 7800 6264 7806 6316
rect 11054 6304 11060 6316
rect 9982 6276 11060 6304
rect 11054 6264 11060 6276
rect 11112 6264 11118 6316
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 11517 6307 11575 6313
rect 11517 6304 11529 6307
rect 11204 6276 11529 6304
rect 11204 6264 11210 6276
rect 11517 6273 11529 6276
rect 11563 6273 11575 6307
rect 13081 6307 13139 6313
rect 13081 6304 13093 6307
rect 11517 6267 11575 6273
rect 11716 6276 13093 6304
rect 2041 6239 2099 6245
rect 2041 6205 2053 6239
rect 2087 6205 2099 6239
rect 2041 6199 2099 6205
rect 6365 6239 6423 6245
rect 6365 6205 6377 6239
rect 6411 6236 6423 6239
rect 8570 6236 8576 6248
rect 6411 6208 8576 6236
rect 6411 6205 6423 6208
rect 6365 6199 6423 6205
rect 2056 6100 2084 6199
rect 8570 6196 8576 6208
rect 8628 6196 8634 6248
rect 8849 6239 8907 6245
rect 8849 6205 8861 6239
rect 8895 6236 8907 6239
rect 8938 6236 8944 6248
rect 8895 6208 8944 6236
rect 8895 6205 8907 6208
rect 8849 6199 8907 6205
rect 8938 6196 8944 6208
rect 8996 6196 9002 6248
rect 10321 6239 10379 6245
rect 10321 6205 10333 6239
rect 10367 6236 10379 6239
rect 11716 6236 11744 6276
rect 13081 6273 13093 6276
rect 13127 6273 13139 6307
rect 13081 6267 13139 6273
rect 13170 6264 13176 6316
rect 13228 6304 13234 6316
rect 13725 6307 13783 6313
rect 13725 6304 13737 6307
rect 13228 6276 13737 6304
rect 13228 6264 13234 6276
rect 13725 6273 13737 6276
rect 13771 6273 13783 6307
rect 13998 6304 14004 6316
rect 13959 6276 14004 6304
rect 13725 6267 13783 6273
rect 13998 6264 14004 6276
rect 14056 6264 14062 6316
rect 14645 6307 14703 6313
rect 14645 6273 14657 6307
rect 14691 6304 14703 6307
rect 15194 6304 15200 6316
rect 14691 6276 15200 6304
rect 14691 6273 14703 6276
rect 14645 6267 14703 6273
rect 15194 6264 15200 6276
rect 15252 6264 15258 6316
rect 12894 6236 12900 6248
rect 10367 6208 11744 6236
rect 12855 6208 12900 6236
rect 10367 6205 10379 6208
rect 10321 6199 10379 6205
rect 12894 6196 12900 6208
rect 12952 6196 12958 6248
rect 13817 6239 13875 6245
rect 13817 6205 13829 6239
rect 13863 6205 13875 6239
rect 13817 6199 13875 6205
rect 13832 6168 13860 6199
rect 10244 6140 13860 6168
rect 2774 6100 2780 6112
rect 2056 6072 2780 6100
rect 2774 6060 2780 6072
rect 2832 6060 2838 6112
rect 3786 6100 3792 6112
rect 3747 6072 3792 6100
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 8662 6060 8668 6112
rect 8720 6100 8726 6112
rect 10244 6100 10272 6140
rect 12802 6100 12808 6112
rect 8720 6072 10272 6100
rect 12763 6072 12808 6100
rect 8720 6060 8726 6072
rect 12802 6060 12808 6072
rect 12860 6060 12866 6112
rect 14001 6103 14059 6109
rect 14001 6069 14013 6103
rect 14047 6100 14059 6103
rect 14550 6100 14556 6112
rect 14047 6072 14556 6100
rect 14047 6069 14059 6072
rect 14001 6063 14059 6069
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 1104 6010 28888 6032
rect 1104 5958 4424 6010
rect 4476 5958 4488 6010
rect 4540 5958 4552 6010
rect 4604 5958 4616 6010
rect 4668 5958 4680 6010
rect 4732 5958 11372 6010
rect 11424 5958 11436 6010
rect 11488 5958 11500 6010
rect 11552 5958 11564 6010
rect 11616 5958 11628 6010
rect 11680 5958 18320 6010
rect 18372 5958 18384 6010
rect 18436 5958 18448 6010
rect 18500 5958 18512 6010
rect 18564 5958 18576 6010
rect 18628 5958 25268 6010
rect 25320 5958 25332 6010
rect 25384 5958 25396 6010
rect 25448 5958 25460 6010
rect 25512 5958 25524 6010
rect 25576 5958 28888 6010
rect 1104 5936 28888 5958
rect 3786 5856 3792 5908
rect 3844 5896 3850 5908
rect 6365 5899 6423 5905
rect 6365 5896 6377 5899
rect 3844 5868 6377 5896
rect 3844 5856 3850 5868
rect 6365 5865 6377 5868
rect 6411 5865 6423 5899
rect 6365 5859 6423 5865
rect 6825 5899 6883 5905
rect 6825 5865 6837 5899
rect 6871 5896 6883 5899
rect 8662 5896 8668 5908
rect 6871 5868 8668 5896
rect 6871 5865 6883 5868
rect 6825 5859 6883 5865
rect 8662 5856 8668 5868
rect 8720 5856 8726 5908
rect 8938 5896 8944 5908
rect 8899 5868 8944 5896
rect 8938 5856 8944 5868
rect 8996 5856 9002 5908
rect 11425 5899 11483 5905
rect 11425 5865 11437 5899
rect 11471 5896 11483 5899
rect 12802 5896 12808 5908
rect 11471 5868 12808 5896
rect 11471 5865 11483 5868
rect 11425 5859 11483 5865
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 11054 5788 11060 5840
rect 11112 5828 11118 5840
rect 13449 5831 13507 5837
rect 13449 5828 13461 5831
rect 11112 5800 13461 5828
rect 11112 5788 11118 5800
rect 13449 5797 13461 5800
rect 13495 5797 13507 5831
rect 13449 5791 13507 5797
rect 6546 5760 6552 5772
rect 6507 5732 6552 5760
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 8570 5720 8576 5772
rect 8628 5760 8634 5772
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 8628 5732 9689 5760
rect 8628 5720 8634 5732
rect 9677 5729 9689 5732
rect 9723 5760 9735 5763
rect 10318 5760 10324 5772
rect 9723 5732 10324 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 10686 5720 10692 5772
rect 10744 5760 10750 5772
rect 16025 5763 16083 5769
rect 16025 5760 16037 5763
rect 10744 5732 16037 5760
rect 10744 5720 10750 5732
rect 16025 5729 16037 5732
rect 16071 5729 16083 5763
rect 16025 5723 16083 5729
rect 6270 5652 6276 5704
rect 6328 5692 6334 5704
rect 6365 5695 6423 5701
rect 6365 5692 6377 5695
rect 6328 5664 6377 5692
rect 6328 5652 6334 5664
rect 6365 5661 6377 5664
rect 6411 5661 6423 5695
rect 6365 5655 6423 5661
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5692 6699 5695
rect 7466 5692 7472 5704
rect 6687 5664 7472 5692
rect 6687 5661 6699 5664
rect 6641 5655 6699 5661
rect 7466 5652 7472 5664
rect 7524 5652 7530 5704
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5661 13599 5695
rect 13541 5655 13599 5661
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5692 14427 5695
rect 15105 5695 15163 5701
rect 15105 5692 15117 5695
rect 14415 5664 15117 5692
rect 14415 5661 14427 5664
rect 14369 5655 14427 5661
rect 15105 5661 15117 5664
rect 15151 5692 15163 5695
rect 15194 5692 15200 5704
rect 15151 5664 15200 5692
rect 15151 5661 15163 5664
rect 15105 5655 15163 5661
rect 9950 5624 9956 5636
rect 9911 5596 9956 5624
rect 9950 5584 9956 5596
rect 10008 5584 10014 5636
rect 13078 5624 13084 5636
rect 11178 5596 13084 5624
rect 13078 5584 13084 5596
rect 13136 5584 13142 5636
rect 13556 5568 13584 5655
rect 15194 5652 15200 5664
rect 15252 5652 15258 5704
rect 15933 5695 15991 5701
rect 15933 5661 15945 5695
rect 15979 5661 15991 5695
rect 15933 5655 15991 5661
rect 15948 5624 15976 5655
rect 14936 5596 15976 5624
rect 13538 5516 13544 5568
rect 13596 5556 13602 5568
rect 14185 5559 14243 5565
rect 14185 5556 14197 5559
rect 13596 5528 14197 5556
rect 13596 5516 13602 5528
rect 14185 5525 14197 5528
rect 14231 5525 14243 5559
rect 14185 5519 14243 5525
rect 14734 5516 14740 5568
rect 14792 5556 14798 5568
rect 14936 5565 14964 5596
rect 14921 5559 14979 5565
rect 14921 5556 14933 5559
rect 14792 5528 14933 5556
rect 14792 5516 14798 5528
rect 14921 5525 14933 5528
rect 14967 5525 14979 5559
rect 14921 5519 14979 5525
rect 1104 5466 28888 5488
rect 1104 5414 7898 5466
rect 7950 5414 7962 5466
rect 8014 5414 8026 5466
rect 8078 5414 8090 5466
rect 8142 5414 8154 5466
rect 8206 5414 14846 5466
rect 14898 5414 14910 5466
rect 14962 5414 14974 5466
rect 15026 5414 15038 5466
rect 15090 5414 15102 5466
rect 15154 5414 21794 5466
rect 21846 5414 21858 5466
rect 21910 5414 21922 5466
rect 21974 5414 21986 5466
rect 22038 5414 22050 5466
rect 22102 5414 28888 5466
rect 1104 5392 28888 5414
rect 8570 5312 8576 5364
rect 8628 5352 8634 5364
rect 9125 5355 9183 5361
rect 9125 5352 9137 5355
rect 8628 5324 9137 5352
rect 8628 5312 8634 5324
rect 9125 5321 9137 5324
rect 9171 5321 9183 5355
rect 9125 5315 9183 5321
rect 4278 5256 6914 5284
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5185 5043 5219
rect 5258 5216 5264 5228
rect 5219 5188 5264 5216
rect 4985 5179 5043 5185
rect 2774 5148 2780 5160
rect 2735 5120 2780 5148
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5148 3111 5151
rect 3786 5148 3792 5160
rect 3099 5120 3792 5148
rect 3099 5117 3111 5120
rect 3053 5111 3111 5117
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5148 4583 5151
rect 5000 5148 5028 5179
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 6886 5216 6914 5256
rect 7650 5244 7656 5296
rect 7708 5284 7714 5296
rect 7837 5287 7895 5293
rect 7837 5284 7849 5287
rect 7708 5256 7849 5284
rect 7708 5244 7714 5256
rect 7837 5253 7849 5256
rect 7883 5253 7895 5287
rect 19886 5284 19892 5296
rect 7837 5247 7895 5253
rect 7944 5256 19892 5284
rect 7944 5216 7972 5256
rect 19886 5244 19892 5256
rect 19944 5244 19950 5296
rect 6886 5188 7972 5216
rect 9950 5176 9956 5228
rect 10008 5216 10014 5228
rect 10045 5219 10103 5225
rect 10045 5216 10057 5219
rect 10008 5188 10057 5216
rect 10008 5176 10014 5188
rect 10045 5185 10057 5188
rect 10091 5185 10103 5219
rect 10045 5179 10103 5185
rect 13817 5219 13875 5225
rect 13817 5185 13829 5219
rect 13863 5216 13875 5219
rect 14274 5216 14280 5228
rect 13863 5188 14280 5216
rect 13863 5185 13875 5188
rect 13817 5179 13875 5185
rect 14274 5176 14280 5188
rect 14332 5216 14338 5228
rect 14642 5216 14648 5228
rect 14332 5188 14648 5216
rect 14332 5176 14338 5188
rect 14642 5176 14648 5188
rect 14700 5176 14706 5228
rect 4571 5120 5028 5148
rect 4571 5117 4583 5120
rect 4525 5111 4583 5117
rect 5074 5108 5080 5160
rect 5132 5148 5138 5160
rect 5132 5120 5177 5148
rect 5132 5108 5138 5120
rect 8110 5108 8116 5160
rect 8168 5148 8174 5160
rect 14090 5148 14096 5160
rect 8168 5120 14096 5148
rect 8168 5108 8174 5120
rect 14090 5108 14096 5120
rect 14148 5108 14154 5160
rect 5445 5083 5503 5089
rect 5445 5049 5457 5083
rect 5491 5080 5503 5083
rect 13170 5080 13176 5092
rect 5491 5052 13176 5080
rect 5491 5049 5503 5052
rect 5445 5043 5503 5049
rect 13170 5040 13176 5052
rect 13228 5040 13234 5092
rect 1762 4972 1768 5024
rect 1820 5012 1826 5024
rect 2133 5015 2191 5021
rect 2133 5012 2145 5015
rect 1820 4984 2145 5012
rect 1820 4972 1826 4984
rect 2133 4981 2145 4984
rect 2179 4981 2191 5015
rect 2133 4975 2191 4981
rect 4890 4972 4896 5024
rect 4948 5012 4954 5024
rect 4985 5015 5043 5021
rect 4985 5012 4997 5015
rect 4948 4984 4997 5012
rect 4948 4972 4954 4984
rect 4985 4981 4997 4984
rect 5031 4981 5043 5015
rect 4985 4975 5043 4981
rect 6638 4972 6644 5024
rect 6696 5012 6702 5024
rect 6733 5015 6791 5021
rect 6733 5012 6745 5015
rect 6696 4984 6745 5012
rect 6696 4972 6702 4984
rect 6733 4981 6745 4984
rect 6779 4981 6791 5015
rect 11698 5012 11704 5024
rect 11659 4984 11704 5012
rect 6733 4975 6791 4981
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 13722 5012 13728 5024
rect 13683 4984 13728 5012
rect 13722 4972 13728 4984
rect 13780 4972 13786 5024
rect 1104 4922 28888 4944
rect 1104 4870 4424 4922
rect 4476 4870 4488 4922
rect 4540 4870 4552 4922
rect 4604 4870 4616 4922
rect 4668 4870 4680 4922
rect 4732 4870 11372 4922
rect 11424 4870 11436 4922
rect 11488 4870 11500 4922
rect 11552 4870 11564 4922
rect 11616 4870 11628 4922
rect 11680 4870 18320 4922
rect 18372 4870 18384 4922
rect 18436 4870 18448 4922
rect 18500 4870 18512 4922
rect 18564 4870 18576 4922
rect 18628 4870 25268 4922
rect 25320 4870 25332 4922
rect 25384 4870 25396 4922
rect 25448 4870 25460 4922
rect 25512 4870 25524 4922
rect 25576 4870 28888 4922
rect 1104 4848 28888 4870
rect 3786 4808 3792 4820
rect 3747 4780 3792 4808
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 8110 4808 8116 4820
rect 8071 4780 8116 4808
rect 8110 4768 8116 4780
rect 8168 4768 8174 4820
rect 13078 4768 13084 4820
rect 13136 4808 13142 4820
rect 13449 4811 13507 4817
rect 13449 4808 13461 4811
rect 13136 4780 13461 4808
rect 13136 4768 13142 4780
rect 13449 4777 13461 4780
rect 13495 4777 13507 4811
rect 13449 4771 13507 4777
rect 14182 4768 14188 4820
rect 14240 4768 14246 4820
rect 16574 4768 16580 4820
rect 16632 4808 16638 4820
rect 16945 4811 17003 4817
rect 16945 4808 16957 4811
rect 16632 4780 16957 4808
rect 16632 4768 16638 4780
rect 16945 4777 16957 4780
rect 16991 4777 17003 4811
rect 19886 4808 19892 4820
rect 19847 4780 19892 4808
rect 16945 4771 17003 4777
rect 19886 4768 19892 4780
rect 19944 4768 19950 4820
rect 3237 4743 3295 4749
rect 3237 4709 3249 4743
rect 3283 4740 3295 4743
rect 5074 4740 5080 4752
rect 3283 4712 5080 4740
rect 3283 4709 3295 4712
rect 3237 4703 3295 4709
rect 5074 4700 5080 4712
rect 5132 4700 5138 4752
rect 12069 4743 12127 4749
rect 12069 4709 12081 4743
rect 12115 4740 12127 4743
rect 14200 4740 14228 4768
rect 12115 4712 14228 4740
rect 12115 4709 12127 4712
rect 12069 4703 12127 4709
rect 1489 4675 1547 4681
rect 1489 4641 1501 4675
rect 1535 4672 1547 4675
rect 2774 4672 2780 4684
rect 1535 4644 2780 4672
rect 1535 4641 1547 4644
rect 1489 4635 1547 4641
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 6362 4672 6368 4684
rect 6323 4644 6368 4672
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 6638 4672 6644 4684
rect 6599 4644 6644 4672
rect 6638 4632 6644 4644
rect 6696 4632 6702 4684
rect 10318 4672 10324 4684
rect 10279 4644 10324 4672
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 10962 4632 10968 4684
rect 11020 4672 11026 4684
rect 14185 4675 14243 4681
rect 14185 4672 14197 4675
rect 11020 4644 14197 4672
rect 11020 4632 11026 4644
rect 14185 4641 14197 4644
rect 14231 4641 14243 4675
rect 14185 4635 14243 4641
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4709 4607 4767 4613
rect 4709 4604 4721 4607
rect 4212 4576 4721 4604
rect 4212 4564 4218 4576
rect 4709 4573 4721 4576
rect 4755 4604 4767 4607
rect 4890 4604 4896 4616
rect 4755 4576 4896 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 4890 4564 4896 4576
rect 4948 4564 4954 4616
rect 13538 4604 13544 4616
rect 13499 4576 13544 4604
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14921 4607 14979 4613
rect 14921 4573 14933 4607
rect 14967 4604 14979 4607
rect 16485 4607 16543 4613
rect 14967 4576 16252 4604
rect 14967 4573 14979 4576
rect 14921 4567 14979 4573
rect 1762 4536 1768 4548
rect 1723 4508 1768 4536
rect 1762 4496 1768 4508
rect 1820 4496 1826 4548
rect 3050 4536 3056 4548
rect 2990 4508 3056 4536
rect 3050 4496 3056 4508
rect 3108 4496 3114 4548
rect 7650 4496 7656 4548
rect 7708 4496 7714 4548
rect 10594 4536 10600 4548
rect 10555 4508 10600 4536
rect 10594 4496 10600 4508
rect 10652 4496 10658 4548
rect 14829 4539 14887 4545
rect 14829 4536 14841 4539
rect 11822 4508 14841 4536
rect 14829 4505 14841 4508
rect 14875 4505 14887 4539
rect 14829 4499 14887 4505
rect 4614 4468 4620 4480
rect 4575 4440 4620 4468
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 13538 4428 13544 4480
rect 13596 4468 13602 4480
rect 14936 4468 14964 4567
rect 16224 4548 16252 4576
rect 16485 4573 16497 4607
rect 16531 4604 16543 4607
rect 16574 4604 16580 4616
rect 16531 4576 16580 4604
rect 16531 4573 16543 4576
rect 16485 4567 16543 4573
rect 16574 4564 16580 4576
rect 16632 4564 16638 4616
rect 19797 4607 19855 4613
rect 19797 4573 19809 4607
rect 19843 4573 19855 4607
rect 19797 4567 19855 4573
rect 16206 4496 16212 4548
rect 16264 4536 16270 4548
rect 19812 4536 19840 4567
rect 16264 4508 19840 4536
rect 16264 4496 16270 4508
rect 16390 4468 16396 4480
rect 13596 4440 14964 4468
rect 16351 4440 16396 4468
rect 13596 4428 13602 4440
rect 16390 4428 16396 4440
rect 16448 4428 16454 4480
rect 1104 4378 28888 4400
rect 1104 4326 7898 4378
rect 7950 4326 7962 4378
rect 8014 4326 8026 4378
rect 8078 4326 8090 4378
rect 8142 4326 8154 4378
rect 8206 4326 14846 4378
rect 14898 4326 14910 4378
rect 14962 4326 14974 4378
rect 15026 4326 15038 4378
rect 15090 4326 15102 4378
rect 15154 4326 21794 4378
rect 21846 4326 21858 4378
rect 21910 4326 21922 4378
rect 21974 4326 21986 4378
rect 22038 4326 22050 4378
rect 22102 4326 28888 4378
rect 1104 4304 28888 4326
rect 16114 4264 16120 4276
rect 11624 4236 16120 4264
rect 4614 4196 4620 4208
rect 3542 4168 4620 4196
rect 4614 4156 4620 4168
rect 4672 4156 4678 4208
rect 11624 4196 11652 4236
rect 16114 4224 16120 4236
rect 16172 4224 16178 4276
rect 7866 4168 11652 4196
rect 11698 4156 11704 4208
rect 11756 4196 11762 4208
rect 11793 4199 11851 4205
rect 11793 4196 11805 4199
rect 11756 4168 11805 4196
rect 11756 4156 11762 4168
rect 11793 4165 11805 4168
rect 11839 4165 11851 4199
rect 13722 4196 13728 4208
rect 13018 4168 13728 4196
rect 11793 4159 11851 4165
rect 13722 4156 13728 4168
rect 13780 4156 13786 4208
rect 6362 4128 6368 4140
rect 6323 4100 6368 4128
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 10318 4088 10324 4140
rect 10376 4128 10382 4140
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 10376 4100 11529 4128
rect 10376 4088 10382 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 2041 4063 2099 4069
rect 2041 4029 2053 4063
rect 2087 4029 2099 4063
rect 2041 4023 2099 4029
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 3050 4060 3056 4072
rect 2363 4032 3056 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 2056 3924 2084 4023
rect 3050 4020 3056 4032
rect 3108 4020 3114 4072
rect 5810 4020 5816 4072
rect 5868 4060 5874 4072
rect 6641 4063 6699 4069
rect 6641 4060 6653 4063
rect 5868 4032 6653 4060
rect 5868 4020 5874 4032
rect 6641 4029 6653 4032
rect 6687 4029 6699 4063
rect 10594 4060 10600 4072
rect 10555 4032 10600 4060
rect 6641 4023 6699 4029
rect 10594 4020 10600 4032
rect 10652 4020 10658 4072
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 14366 4060 14372 4072
rect 13311 4032 14372 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 2774 3924 2780 3936
rect 2056 3896 2780 3924
rect 2774 3884 2780 3896
rect 2832 3884 2838 3936
rect 3789 3927 3847 3933
rect 3789 3893 3801 3927
rect 3835 3924 3847 3927
rect 8018 3924 8024 3936
rect 3835 3896 8024 3924
rect 3835 3893 3847 3896
rect 3789 3887 3847 3893
rect 8018 3884 8024 3896
rect 8076 3884 8082 3936
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3924 8171 3927
rect 12894 3924 12900 3936
rect 8159 3896 12900 3924
rect 8159 3893 8171 3896
rect 8113 3887 8171 3893
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 1104 3834 28888 3856
rect 1104 3782 4424 3834
rect 4476 3782 4488 3834
rect 4540 3782 4552 3834
rect 4604 3782 4616 3834
rect 4668 3782 4680 3834
rect 4732 3782 11372 3834
rect 11424 3782 11436 3834
rect 11488 3782 11500 3834
rect 11552 3782 11564 3834
rect 11616 3782 11628 3834
rect 11680 3782 18320 3834
rect 18372 3782 18384 3834
rect 18436 3782 18448 3834
rect 18500 3782 18512 3834
rect 18564 3782 18576 3834
rect 18628 3782 25268 3834
rect 25320 3782 25332 3834
rect 25384 3782 25396 3834
rect 25448 3782 25460 3834
rect 25512 3782 25524 3834
rect 25576 3782 28888 3834
rect 1104 3760 28888 3782
rect 14 3680 20 3732
rect 72 3720 78 3732
rect 6086 3720 6092 3732
rect 72 3692 6092 3720
rect 72 3680 78 3692
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 12161 3723 12219 3729
rect 6288 3692 10548 3720
rect 3050 3652 3056 3664
rect 3011 3624 3056 3652
rect 3050 3612 3056 3624
rect 3108 3612 3114 3664
rect 5721 3655 5779 3661
rect 5721 3621 5733 3655
rect 5767 3652 5779 3655
rect 6288 3652 6316 3692
rect 5767 3624 6316 3652
rect 5767 3621 5779 3624
rect 5721 3615 5779 3621
rect 7466 3612 7472 3664
rect 7524 3652 7530 3664
rect 7929 3655 7987 3661
rect 7929 3652 7941 3655
rect 7524 3624 7941 3652
rect 7524 3612 7530 3624
rect 7929 3621 7941 3624
rect 7975 3621 7987 3655
rect 7929 3615 7987 3621
rect 2774 3544 2780 3596
rect 2832 3584 2838 3596
rect 3973 3587 4031 3593
rect 3973 3584 3985 3587
rect 2832 3556 3985 3584
rect 2832 3544 2838 3556
rect 3973 3553 3985 3556
rect 4019 3584 4031 3587
rect 4019 3556 6224 3584
rect 4019 3553 4031 3556
rect 3973 3547 4031 3553
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3485 2007 3519
rect 1949 3479 2007 3485
rect 1964 3448 1992 3479
rect 2038 3476 2044 3528
rect 2096 3516 2102 3528
rect 6196 3525 6224 3556
rect 10318 3544 10324 3596
rect 10376 3584 10382 3596
rect 10413 3587 10471 3593
rect 10413 3584 10425 3587
rect 10376 3556 10425 3584
rect 10376 3544 10382 3556
rect 10413 3553 10425 3556
rect 10459 3553 10471 3587
rect 10520 3584 10548 3692
rect 12161 3689 12173 3723
rect 12207 3720 12219 3723
rect 14645 3723 14703 3729
rect 14645 3720 14657 3723
rect 12207 3692 14657 3720
rect 12207 3689 12219 3692
rect 12161 3683 12219 3689
rect 14645 3689 14657 3692
rect 14691 3689 14703 3723
rect 16114 3720 16120 3732
rect 16075 3692 16120 3720
rect 14645 3683 14703 3689
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 13998 3612 14004 3664
rect 14056 3652 14062 3664
rect 15105 3655 15163 3661
rect 15105 3652 15117 3655
rect 14056 3624 15117 3652
rect 14056 3612 14062 3624
rect 15105 3621 15117 3624
rect 15151 3621 15163 3655
rect 15105 3615 15163 3621
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 10520 3556 14749 3584
rect 10413 3547 10471 3553
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 2409 3519 2467 3525
rect 2409 3516 2421 3519
rect 2096 3488 2421 3516
rect 2096 3476 2102 3488
rect 2409 3485 2421 3488
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3485 6239 3519
rect 6181 3479 6239 3485
rect 3970 3448 3976 3460
rect 1964 3420 3976 3448
rect 3970 3408 3976 3420
rect 4028 3408 4034 3460
rect 4246 3448 4252 3460
rect 4207 3420 4252 3448
rect 4246 3408 4252 3420
rect 4304 3408 4310 3460
rect 6196 3448 6224 3479
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8536 3488 8953 3516
rect 8536 3476 8542 3488
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 11974 3476 11980 3528
rect 12032 3516 12038 3528
rect 14921 3519 14979 3525
rect 14921 3516 14933 3519
rect 12032 3488 14933 3516
rect 12032 3476 12038 3488
rect 14921 3485 14933 3488
rect 14967 3485 14979 3519
rect 16206 3516 16212 3528
rect 16167 3488 16212 3516
rect 14921 3479 14979 3485
rect 16206 3476 16212 3488
rect 16264 3476 16270 3528
rect 6362 3448 6368 3460
rect 4356 3420 4738 3448
rect 6196 3420 6368 3448
rect 1857 3383 1915 3389
rect 1857 3349 1869 3383
rect 1903 3380 1915 3383
rect 4356 3380 4384 3420
rect 6362 3408 6368 3420
rect 6420 3408 6426 3460
rect 6457 3451 6515 3457
rect 6457 3417 6469 3451
rect 6503 3448 6515 3451
rect 6546 3448 6552 3460
rect 6503 3420 6552 3448
rect 6503 3417 6515 3420
rect 6457 3411 6515 3417
rect 6546 3408 6552 3420
rect 6604 3408 6610 3460
rect 10594 3448 10600 3460
rect 7682 3420 10600 3448
rect 10594 3408 10600 3420
rect 10652 3408 10658 3460
rect 10689 3451 10747 3457
rect 10689 3417 10701 3451
rect 10735 3448 10747 3451
rect 10778 3448 10784 3460
rect 10735 3420 10784 3448
rect 10735 3417 10747 3420
rect 10689 3411 10747 3417
rect 10778 3408 10784 3420
rect 10836 3408 10842 3460
rect 14458 3448 14464 3460
rect 11914 3420 14464 3448
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 14645 3451 14703 3457
rect 14645 3417 14657 3451
rect 14691 3417 14703 3451
rect 14645 3411 14703 3417
rect 1903 3352 4384 3380
rect 1903 3349 1915 3352
rect 1857 3343 1915 3349
rect 4890 3340 4896 3392
rect 4948 3380 4954 3392
rect 7742 3380 7748 3392
rect 4948 3352 7748 3380
rect 4948 3340 4954 3352
rect 7742 3340 7748 3352
rect 7800 3340 7806 3392
rect 8018 3340 8024 3392
rect 8076 3380 8082 3392
rect 14660 3380 14688 3411
rect 8076 3352 14688 3380
rect 8076 3340 8082 3352
rect 1104 3290 28888 3312
rect 1104 3238 7898 3290
rect 7950 3238 7962 3290
rect 8014 3238 8026 3290
rect 8078 3238 8090 3290
rect 8142 3238 8154 3290
rect 8206 3238 14846 3290
rect 14898 3238 14910 3290
rect 14962 3238 14974 3290
rect 15026 3238 15038 3290
rect 15090 3238 15102 3290
rect 15154 3238 21794 3290
rect 21846 3238 21858 3290
rect 21910 3238 21922 3290
rect 21974 3238 21986 3290
rect 22038 3238 22050 3290
rect 22102 3238 28888 3290
rect 1104 3216 28888 3238
rect 10318 3176 10324 3188
rect 8220 3148 10324 3176
rect 2774 3108 2780 3120
rect 2735 3080 2780 3108
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 4338 3108 4344 3120
rect 4299 3080 4344 3108
rect 4338 3068 4344 3080
rect 4396 3068 4402 3120
rect 4246 3000 4252 3052
rect 4304 3040 4310 3052
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4304 3012 4997 3040
rect 4304 3000 4310 3012
rect 4985 3009 4997 3012
rect 5031 3009 5043 3043
rect 5810 3040 5816 3052
rect 5771 3012 5816 3040
rect 4985 3003 5043 3009
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 6546 3040 6552 3052
rect 6507 3012 6552 3040
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 8220 3049 8248 3148
rect 10318 3136 10324 3148
rect 10376 3136 10382 3188
rect 10594 3136 10600 3188
rect 10652 3176 10658 3188
rect 14458 3176 14464 3188
rect 10652 3148 11100 3176
rect 14419 3148 14464 3176
rect 10652 3136 10658 3148
rect 8478 3108 8484 3120
rect 8439 3080 8484 3108
rect 8478 3068 8484 3080
rect 8536 3068 8542 3120
rect 10962 3108 10968 3120
rect 9706 3080 10968 3108
rect 10962 3068 10968 3080
rect 11020 3068 11026 3120
rect 11072 3108 11100 3148
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 15105 3111 15163 3117
rect 15105 3108 15117 3111
rect 11072 3080 15117 3108
rect 15105 3077 15117 3080
rect 15151 3077 15163 3111
rect 15105 3071 15163 3077
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3009 8263 3043
rect 10778 3040 10784 3052
rect 10739 3012 10784 3040
rect 8205 3003 8263 3009
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3040 14611 3043
rect 14734 3040 14740 3052
rect 14599 3012 14740 3040
rect 14599 3009 14611 3012
rect 14553 3003 14611 3009
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 9953 2975 10011 2981
rect 7800 2944 9904 2972
rect 7800 2932 7806 2944
rect 9876 2904 9904 2944
rect 9953 2941 9965 2975
rect 9999 2972 10011 2975
rect 11974 2972 11980 2984
rect 9999 2944 11980 2972
rect 9999 2941 10011 2944
rect 9953 2935 10011 2941
rect 11974 2932 11980 2944
rect 12032 2932 12038 2984
rect 14568 2904 14596 3003
rect 14734 3000 14740 3012
rect 14792 3040 14798 3052
rect 15197 3043 15255 3049
rect 15197 3040 15209 3043
rect 14792 3012 15209 3040
rect 14792 3000 14798 3012
rect 15197 3009 15209 3012
rect 15243 3009 15255 3043
rect 15197 3003 15255 3009
rect 9876 2876 14596 2904
rect 1104 2746 28888 2768
rect 1104 2694 4424 2746
rect 4476 2694 4488 2746
rect 4540 2694 4552 2746
rect 4604 2694 4616 2746
rect 4668 2694 4680 2746
rect 4732 2694 11372 2746
rect 11424 2694 11436 2746
rect 11488 2694 11500 2746
rect 11552 2694 11564 2746
rect 11616 2694 11628 2746
rect 11680 2694 18320 2746
rect 18372 2694 18384 2746
rect 18436 2694 18448 2746
rect 18500 2694 18512 2746
rect 18564 2694 18576 2746
rect 18628 2694 25268 2746
rect 25320 2694 25332 2746
rect 25384 2694 25396 2746
rect 25448 2694 25460 2746
rect 25512 2694 25524 2746
rect 25576 2694 28888 2746
rect 1104 2672 28888 2694
rect 3237 2635 3295 2641
rect 3237 2601 3249 2635
rect 3283 2632 3295 2635
rect 5258 2632 5264 2644
rect 3283 2604 5264 2632
rect 3283 2601 3295 2604
rect 3237 2595 3295 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 23290 2564 23296 2576
rect 23251 2536 23296 2564
rect 23290 2524 23296 2536
rect 23348 2524 23354 2576
rect 1489 2499 1547 2505
rect 1489 2465 1501 2499
rect 1535 2496 1547 2499
rect 2774 2496 2780 2508
rect 1535 2468 2780 2496
rect 1535 2465 1547 2468
rect 1489 2459 1547 2465
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 1765 2363 1823 2369
rect 1765 2329 1777 2363
rect 1811 2360 1823 2363
rect 2038 2360 2044 2372
rect 1811 2332 2044 2360
rect 1811 2329 1823 2332
rect 1765 2323 1823 2329
rect 2038 2320 2044 2332
rect 2096 2320 2102 2372
rect 16390 2360 16396 2372
rect 2990 2332 16396 2360
rect 16390 2320 16396 2332
rect 16448 2320 16454 2372
rect 22833 2363 22891 2369
rect 22833 2329 22845 2363
rect 22879 2360 22891 2363
rect 23198 2360 23204 2372
rect 22879 2332 23204 2360
rect 22879 2329 22891 2332
rect 22833 2323 22891 2329
rect 23198 2320 23204 2332
rect 23256 2360 23262 2372
rect 23477 2363 23535 2369
rect 23477 2360 23489 2363
rect 23256 2332 23489 2360
rect 23256 2320 23262 2332
rect 23477 2329 23489 2332
rect 23523 2329 23535 2363
rect 23477 2323 23535 2329
rect 1104 2202 28888 2224
rect 1104 2150 7898 2202
rect 7950 2150 7962 2202
rect 8014 2150 8026 2202
rect 8078 2150 8090 2202
rect 8142 2150 8154 2202
rect 8206 2150 14846 2202
rect 14898 2150 14910 2202
rect 14962 2150 14974 2202
rect 15026 2150 15038 2202
rect 15090 2150 15102 2202
rect 15154 2150 21794 2202
rect 21846 2150 21858 2202
rect 21910 2150 21922 2202
rect 21974 2150 21986 2202
rect 22038 2150 22050 2202
rect 22102 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 4424 27718 4476 27770
rect 4488 27718 4540 27770
rect 4552 27718 4604 27770
rect 4616 27718 4668 27770
rect 4680 27718 4732 27770
rect 11372 27718 11424 27770
rect 11436 27718 11488 27770
rect 11500 27718 11552 27770
rect 11564 27718 11616 27770
rect 11628 27718 11680 27770
rect 18320 27718 18372 27770
rect 18384 27718 18436 27770
rect 18448 27718 18500 27770
rect 18512 27718 18564 27770
rect 18576 27718 18628 27770
rect 25268 27718 25320 27770
rect 25332 27718 25384 27770
rect 25396 27718 25448 27770
rect 25460 27718 25512 27770
rect 25524 27718 25576 27770
rect 18052 27548 18104 27600
rect 18144 27319 18196 27328
rect 18144 27285 18153 27319
rect 18153 27285 18187 27319
rect 18187 27285 18196 27319
rect 18144 27276 18196 27285
rect 7898 27174 7950 27226
rect 7962 27174 8014 27226
rect 8026 27174 8078 27226
rect 8090 27174 8142 27226
rect 8154 27174 8206 27226
rect 14846 27174 14898 27226
rect 14910 27174 14962 27226
rect 14974 27174 15026 27226
rect 15038 27174 15090 27226
rect 15102 27174 15154 27226
rect 21794 27174 21846 27226
rect 21858 27174 21910 27226
rect 21922 27174 21974 27226
rect 21986 27174 22038 27226
rect 22050 27174 22102 27226
rect 4424 26630 4476 26682
rect 4488 26630 4540 26682
rect 4552 26630 4604 26682
rect 4616 26630 4668 26682
rect 4680 26630 4732 26682
rect 11372 26630 11424 26682
rect 11436 26630 11488 26682
rect 11500 26630 11552 26682
rect 11564 26630 11616 26682
rect 11628 26630 11680 26682
rect 18320 26630 18372 26682
rect 18384 26630 18436 26682
rect 18448 26630 18500 26682
rect 18512 26630 18564 26682
rect 18576 26630 18628 26682
rect 25268 26630 25320 26682
rect 25332 26630 25384 26682
rect 25396 26630 25448 26682
rect 25460 26630 25512 26682
rect 25524 26630 25576 26682
rect 7898 26086 7950 26138
rect 7962 26086 8014 26138
rect 8026 26086 8078 26138
rect 8090 26086 8142 26138
rect 8154 26086 8206 26138
rect 14846 26086 14898 26138
rect 14910 26086 14962 26138
rect 14974 26086 15026 26138
rect 15038 26086 15090 26138
rect 15102 26086 15154 26138
rect 21794 26086 21846 26138
rect 21858 26086 21910 26138
rect 21922 26086 21974 26138
rect 21986 26086 22038 26138
rect 22050 26086 22102 26138
rect 4424 25542 4476 25594
rect 4488 25542 4540 25594
rect 4552 25542 4604 25594
rect 4616 25542 4668 25594
rect 4680 25542 4732 25594
rect 11372 25542 11424 25594
rect 11436 25542 11488 25594
rect 11500 25542 11552 25594
rect 11564 25542 11616 25594
rect 11628 25542 11680 25594
rect 18320 25542 18372 25594
rect 18384 25542 18436 25594
rect 18448 25542 18500 25594
rect 18512 25542 18564 25594
rect 18576 25542 18628 25594
rect 25268 25542 25320 25594
rect 25332 25542 25384 25594
rect 25396 25542 25448 25594
rect 25460 25542 25512 25594
rect 25524 25542 25576 25594
rect 7898 24998 7950 25050
rect 7962 24998 8014 25050
rect 8026 24998 8078 25050
rect 8090 24998 8142 25050
rect 8154 24998 8206 25050
rect 14846 24998 14898 25050
rect 14910 24998 14962 25050
rect 14974 24998 15026 25050
rect 15038 24998 15090 25050
rect 15102 24998 15154 25050
rect 21794 24998 21846 25050
rect 21858 24998 21910 25050
rect 21922 24998 21974 25050
rect 21986 24998 22038 25050
rect 22050 24998 22102 25050
rect 6368 24760 6420 24812
rect 1492 24599 1544 24608
rect 1492 24565 1501 24599
rect 1501 24565 1535 24599
rect 1535 24565 1544 24599
rect 1492 24556 1544 24565
rect 4424 24454 4476 24506
rect 4488 24454 4540 24506
rect 4552 24454 4604 24506
rect 4616 24454 4668 24506
rect 4680 24454 4732 24506
rect 11372 24454 11424 24506
rect 11436 24454 11488 24506
rect 11500 24454 11552 24506
rect 11564 24454 11616 24506
rect 11628 24454 11680 24506
rect 18320 24454 18372 24506
rect 18384 24454 18436 24506
rect 18448 24454 18500 24506
rect 18512 24454 18564 24506
rect 18576 24454 18628 24506
rect 25268 24454 25320 24506
rect 25332 24454 25384 24506
rect 25396 24454 25448 24506
rect 25460 24454 25512 24506
rect 25524 24454 25576 24506
rect 7898 23910 7950 23962
rect 7962 23910 8014 23962
rect 8026 23910 8078 23962
rect 8090 23910 8142 23962
rect 8154 23910 8206 23962
rect 14846 23910 14898 23962
rect 14910 23910 14962 23962
rect 14974 23910 15026 23962
rect 15038 23910 15090 23962
rect 15102 23910 15154 23962
rect 21794 23910 21846 23962
rect 21858 23910 21910 23962
rect 21922 23910 21974 23962
rect 21986 23910 22038 23962
rect 22050 23910 22102 23962
rect 4424 23366 4476 23418
rect 4488 23366 4540 23418
rect 4552 23366 4604 23418
rect 4616 23366 4668 23418
rect 4680 23366 4732 23418
rect 11372 23366 11424 23418
rect 11436 23366 11488 23418
rect 11500 23366 11552 23418
rect 11564 23366 11616 23418
rect 11628 23366 11680 23418
rect 18320 23366 18372 23418
rect 18384 23366 18436 23418
rect 18448 23366 18500 23418
rect 18512 23366 18564 23418
rect 18576 23366 18628 23418
rect 25268 23366 25320 23418
rect 25332 23366 25384 23418
rect 25396 23366 25448 23418
rect 25460 23366 25512 23418
rect 25524 23366 25576 23418
rect 7898 22822 7950 22874
rect 7962 22822 8014 22874
rect 8026 22822 8078 22874
rect 8090 22822 8142 22874
rect 8154 22822 8206 22874
rect 14846 22822 14898 22874
rect 14910 22822 14962 22874
rect 14974 22822 15026 22874
rect 15038 22822 15090 22874
rect 15102 22822 15154 22874
rect 21794 22822 21846 22874
rect 21858 22822 21910 22874
rect 21922 22822 21974 22874
rect 21986 22822 22038 22874
rect 22050 22822 22102 22874
rect 4424 22278 4476 22330
rect 4488 22278 4540 22330
rect 4552 22278 4604 22330
rect 4616 22278 4668 22330
rect 4680 22278 4732 22330
rect 11372 22278 11424 22330
rect 11436 22278 11488 22330
rect 11500 22278 11552 22330
rect 11564 22278 11616 22330
rect 11628 22278 11680 22330
rect 18320 22278 18372 22330
rect 18384 22278 18436 22330
rect 18448 22278 18500 22330
rect 18512 22278 18564 22330
rect 18576 22278 18628 22330
rect 25268 22278 25320 22330
rect 25332 22278 25384 22330
rect 25396 22278 25448 22330
rect 25460 22278 25512 22330
rect 25524 22278 25576 22330
rect 7898 21734 7950 21786
rect 7962 21734 8014 21786
rect 8026 21734 8078 21786
rect 8090 21734 8142 21786
rect 8154 21734 8206 21786
rect 14846 21734 14898 21786
rect 14910 21734 14962 21786
rect 14974 21734 15026 21786
rect 15038 21734 15090 21786
rect 15102 21734 15154 21786
rect 21794 21734 21846 21786
rect 21858 21734 21910 21786
rect 21922 21734 21974 21786
rect 21986 21734 22038 21786
rect 22050 21734 22102 21786
rect 4424 21190 4476 21242
rect 4488 21190 4540 21242
rect 4552 21190 4604 21242
rect 4616 21190 4668 21242
rect 4680 21190 4732 21242
rect 11372 21190 11424 21242
rect 11436 21190 11488 21242
rect 11500 21190 11552 21242
rect 11564 21190 11616 21242
rect 11628 21190 11680 21242
rect 18320 21190 18372 21242
rect 18384 21190 18436 21242
rect 18448 21190 18500 21242
rect 18512 21190 18564 21242
rect 18576 21190 18628 21242
rect 25268 21190 25320 21242
rect 25332 21190 25384 21242
rect 25396 21190 25448 21242
rect 25460 21190 25512 21242
rect 25524 21190 25576 21242
rect 7898 20646 7950 20698
rect 7962 20646 8014 20698
rect 8026 20646 8078 20698
rect 8090 20646 8142 20698
rect 8154 20646 8206 20698
rect 14846 20646 14898 20698
rect 14910 20646 14962 20698
rect 14974 20646 15026 20698
rect 15038 20646 15090 20698
rect 15102 20646 15154 20698
rect 21794 20646 21846 20698
rect 21858 20646 21910 20698
rect 21922 20646 21974 20698
rect 21986 20646 22038 20698
rect 22050 20646 22102 20698
rect 3976 20408 4028 20460
rect 3792 20204 3844 20256
rect 3976 20247 4028 20256
rect 3976 20213 3985 20247
rect 3985 20213 4019 20247
rect 4019 20213 4028 20247
rect 3976 20204 4028 20213
rect 4424 20102 4476 20154
rect 4488 20102 4540 20154
rect 4552 20102 4604 20154
rect 4616 20102 4668 20154
rect 4680 20102 4732 20154
rect 11372 20102 11424 20154
rect 11436 20102 11488 20154
rect 11500 20102 11552 20154
rect 11564 20102 11616 20154
rect 11628 20102 11680 20154
rect 18320 20102 18372 20154
rect 18384 20102 18436 20154
rect 18448 20102 18500 20154
rect 18512 20102 18564 20154
rect 18576 20102 18628 20154
rect 25268 20102 25320 20154
rect 25332 20102 25384 20154
rect 25396 20102 25448 20154
rect 25460 20102 25512 20154
rect 25524 20102 25576 20154
rect 3148 19796 3200 19848
rect 3976 19796 4028 19848
rect 3424 19660 3476 19712
rect 7898 19558 7950 19610
rect 7962 19558 8014 19610
rect 8026 19558 8078 19610
rect 8090 19558 8142 19610
rect 8154 19558 8206 19610
rect 14846 19558 14898 19610
rect 14910 19558 14962 19610
rect 14974 19558 15026 19610
rect 15038 19558 15090 19610
rect 15102 19558 15154 19610
rect 21794 19558 21846 19610
rect 21858 19558 21910 19610
rect 21922 19558 21974 19610
rect 21986 19558 22038 19610
rect 22050 19558 22102 19610
rect 4424 19014 4476 19066
rect 4488 19014 4540 19066
rect 4552 19014 4604 19066
rect 4616 19014 4668 19066
rect 4680 19014 4732 19066
rect 11372 19014 11424 19066
rect 11436 19014 11488 19066
rect 11500 19014 11552 19066
rect 11564 19014 11616 19066
rect 11628 19014 11680 19066
rect 18320 19014 18372 19066
rect 18384 19014 18436 19066
rect 18448 19014 18500 19066
rect 18512 19014 18564 19066
rect 18576 19014 18628 19066
rect 25268 19014 25320 19066
rect 25332 19014 25384 19066
rect 25396 19014 25448 19066
rect 25460 19014 25512 19066
rect 25524 19014 25576 19066
rect 7898 18470 7950 18522
rect 7962 18470 8014 18522
rect 8026 18470 8078 18522
rect 8090 18470 8142 18522
rect 8154 18470 8206 18522
rect 14846 18470 14898 18522
rect 14910 18470 14962 18522
rect 14974 18470 15026 18522
rect 15038 18470 15090 18522
rect 15102 18470 15154 18522
rect 21794 18470 21846 18522
rect 21858 18470 21910 18522
rect 21922 18470 21974 18522
rect 21986 18470 22038 18522
rect 22050 18470 22102 18522
rect 4424 17926 4476 17978
rect 4488 17926 4540 17978
rect 4552 17926 4604 17978
rect 4616 17926 4668 17978
rect 4680 17926 4732 17978
rect 11372 17926 11424 17978
rect 11436 17926 11488 17978
rect 11500 17926 11552 17978
rect 11564 17926 11616 17978
rect 11628 17926 11680 17978
rect 18320 17926 18372 17978
rect 18384 17926 18436 17978
rect 18448 17926 18500 17978
rect 18512 17926 18564 17978
rect 18576 17926 18628 17978
rect 25268 17926 25320 17978
rect 25332 17926 25384 17978
rect 25396 17926 25448 17978
rect 25460 17926 25512 17978
rect 25524 17926 25576 17978
rect 7898 17382 7950 17434
rect 7962 17382 8014 17434
rect 8026 17382 8078 17434
rect 8090 17382 8142 17434
rect 8154 17382 8206 17434
rect 14846 17382 14898 17434
rect 14910 17382 14962 17434
rect 14974 17382 15026 17434
rect 15038 17382 15090 17434
rect 15102 17382 15154 17434
rect 21794 17382 21846 17434
rect 21858 17382 21910 17434
rect 21922 17382 21974 17434
rect 21986 17382 22038 17434
rect 22050 17382 22102 17434
rect 5632 17212 5684 17264
rect 7564 17212 7616 17264
rect 4896 17144 4948 17196
rect 28172 17187 28224 17196
rect 4988 17008 5040 17060
rect 7380 17008 7432 17060
rect 28172 17153 28181 17187
rect 28181 17153 28215 17187
rect 28215 17153 28224 17187
rect 28172 17144 28224 17153
rect 7932 17119 7984 17128
rect 7932 17085 7941 17119
rect 7941 17085 7975 17119
rect 7975 17085 7984 17119
rect 9036 17119 9088 17128
rect 7932 17076 7984 17085
rect 9036 17085 9045 17119
rect 9045 17085 9079 17119
rect 9079 17085 9088 17119
rect 9036 17076 9088 17085
rect 10324 17076 10376 17128
rect 4804 16940 4856 16992
rect 7656 16940 7708 16992
rect 10416 16940 10468 16992
rect 27988 16983 28040 16992
rect 27988 16949 27997 16983
rect 27997 16949 28031 16983
rect 28031 16949 28040 16983
rect 27988 16940 28040 16949
rect 4424 16838 4476 16890
rect 4488 16838 4540 16890
rect 4552 16838 4604 16890
rect 4616 16838 4668 16890
rect 4680 16838 4732 16890
rect 11372 16838 11424 16890
rect 11436 16838 11488 16890
rect 11500 16838 11552 16890
rect 11564 16838 11616 16890
rect 11628 16838 11680 16890
rect 18320 16838 18372 16890
rect 18384 16838 18436 16890
rect 18448 16838 18500 16890
rect 18512 16838 18564 16890
rect 18576 16838 18628 16890
rect 25268 16838 25320 16890
rect 25332 16838 25384 16890
rect 25396 16838 25448 16890
rect 25460 16838 25512 16890
rect 25524 16838 25576 16890
rect 7932 16736 7984 16788
rect 5632 16600 5684 16652
rect 4804 16575 4856 16584
rect 4804 16541 4813 16575
rect 4813 16541 4847 16575
rect 4847 16541 4856 16575
rect 4804 16532 4856 16541
rect 4988 16575 5040 16584
rect 4988 16541 4997 16575
rect 4997 16541 5031 16575
rect 5031 16541 5040 16575
rect 4988 16532 5040 16541
rect 2964 16464 3016 16516
rect 5724 16532 5776 16584
rect 7564 16600 7616 16652
rect 7748 16643 7800 16652
rect 7748 16609 7757 16643
rect 7757 16609 7791 16643
rect 7791 16609 7800 16643
rect 7748 16600 7800 16609
rect 10416 16668 10468 16720
rect 9312 16575 9364 16584
rect 4068 16396 4120 16448
rect 6644 16464 6696 16516
rect 9312 16541 9321 16575
rect 9321 16541 9355 16575
rect 9355 16541 9364 16575
rect 9312 16532 9364 16541
rect 9588 16575 9640 16584
rect 9588 16541 9597 16575
rect 9597 16541 9631 16575
rect 9631 16541 9640 16575
rect 9588 16532 9640 16541
rect 10324 16575 10376 16584
rect 10324 16541 10333 16575
rect 10333 16541 10367 16575
rect 10367 16541 10376 16575
rect 10324 16532 10376 16541
rect 11704 16532 11756 16584
rect 12440 16532 12492 16584
rect 5540 16439 5592 16448
rect 5540 16405 5549 16439
rect 5549 16405 5583 16439
rect 5583 16405 5592 16439
rect 5540 16396 5592 16405
rect 5724 16396 5776 16448
rect 9588 16396 9640 16448
rect 11704 16439 11756 16448
rect 11704 16405 11713 16439
rect 11713 16405 11747 16439
rect 11747 16405 11756 16439
rect 11704 16396 11756 16405
rect 7898 16294 7950 16346
rect 7962 16294 8014 16346
rect 8026 16294 8078 16346
rect 8090 16294 8142 16346
rect 8154 16294 8206 16346
rect 14846 16294 14898 16346
rect 14910 16294 14962 16346
rect 14974 16294 15026 16346
rect 15038 16294 15090 16346
rect 15102 16294 15154 16346
rect 21794 16294 21846 16346
rect 21858 16294 21910 16346
rect 21922 16294 21974 16346
rect 21986 16294 22038 16346
rect 22050 16294 22102 16346
rect 4896 16192 4948 16244
rect 7748 16192 7800 16244
rect 9312 16235 9364 16244
rect 9312 16201 9321 16235
rect 9321 16201 9355 16235
rect 9355 16201 9364 16235
rect 9312 16192 9364 16201
rect 5540 16124 5592 16176
rect 4896 16099 4948 16108
rect 4896 16065 4905 16099
rect 4905 16065 4939 16099
rect 4939 16065 4948 16099
rect 4896 16056 4948 16065
rect 4988 16099 5040 16108
rect 4988 16065 4997 16099
rect 4997 16065 5031 16099
rect 5031 16065 5040 16099
rect 4988 16056 5040 16065
rect 5448 16056 5500 16108
rect 5724 16056 5776 16108
rect 6644 16099 6696 16108
rect 6644 16065 6653 16099
rect 6653 16065 6687 16099
rect 6687 16065 6696 16099
rect 6644 16056 6696 16065
rect 7380 16056 7432 16108
rect 12440 16056 12492 16108
rect 12992 16056 13044 16108
rect 3792 15988 3844 16040
rect 4160 15988 4212 16040
rect 7472 15988 7524 16040
rect 7656 15988 7708 16040
rect 8300 15988 8352 16040
rect 9036 16031 9088 16040
rect 9036 15997 9045 16031
rect 9045 15997 9079 16031
rect 9079 15997 9088 16031
rect 9036 15988 9088 15997
rect 9404 15988 9456 16040
rect 6368 15963 6420 15972
rect 6368 15929 6377 15963
rect 6377 15929 6411 15963
rect 6411 15929 6420 15963
rect 6368 15920 6420 15929
rect 7196 15852 7248 15904
rect 11796 15895 11848 15904
rect 11796 15861 11805 15895
rect 11805 15861 11839 15895
rect 11839 15861 11848 15895
rect 11796 15852 11848 15861
rect 12164 15895 12216 15904
rect 12164 15861 12173 15895
rect 12173 15861 12207 15895
rect 12207 15861 12216 15895
rect 12164 15852 12216 15861
rect 4424 15750 4476 15802
rect 4488 15750 4540 15802
rect 4552 15750 4604 15802
rect 4616 15750 4668 15802
rect 4680 15750 4732 15802
rect 11372 15750 11424 15802
rect 11436 15750 11488 15802
rect 11500 15750 11552 15802
rect 11564 15750 11616 15802
rect 11628 15750 11680 15802
rect 18320 15750 18372 15802
rect 18384 15750 18436 15802
rect 18448 15750 18500 15802
rect 18512 15750 18564 15802
rect 18576 15750 18628 15802
rect 25268 15750 25320 15802
rect 25332 15750 25384 15802
rect 25396 15750 25448 15802
rect 25460 15750 25512 15802
rect 25524 15750 25576 15802
rect 5632 15648 5684 15700
rect 7380 15691 7432 15700
rect 7380 15657 7389 15691
rect 7389 15657 7423 15691
rect 7423 15657 7432 15691
rect 7380 15648 7432 15657
rect 11704 15648 11756 15700
rect 4988 15512 5040 15564
rect 9864 15580 9916 15632
rect 6736 15512 6788 15564
rect 9496 15512 9548 15564
rect 5724 15487 5776 15496
rect 5724 15453 5733 15487
rect 5733 15453 5767 15487
rect 5767 15453 5776 15487
rect 5724 15444 5776 15453
rect 6368 15444 6420 15496
rect 6644 15487 6696 15496
rect 6644 15453 6653 15487
rect 6653 15453 6687 15487
rect 6687 15453 6696 15487
rect 6644 15444 6696 15453
rect 7380 15444 7432 15496
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 9312 15487 9364 15496
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 9404 15487 9456 15496
rect 9404 15453 9413 15487
rect 9413 15453 9447 15487
rect 9447 15453 9456 15487
rect 9404 15444 9456 15453
rect 11152 15444 11204 15496
rect 14280 15580 14332 15632
rect 5448 15351 5500 15360
rect 5448 15317 5457 15351
rect 5457 15317 5491 15351
rect 5491 15317 5500 15351
rect 5448 15308 5500 15317
rect 5632 15351 5684 15360
rect 5632 15317 5641 15351
rect 5641 15317 5675 15351
rect 5675 15317 5684 15351
rect 5632 15308 5684 15317
rect 8300 15308 8352 15360
rect 8760 15308 8812 15360
rect 11888 15351 11940 15360
rect 11888 15317 11897 15351
rect 11897 15317 11931 15351
rect 11931 15317 11940 15351
rect 11888 15308 11940 15317
rect 12808 15351 12860 15360
rect 12808 15317 12817 15351
rect 12817 15317 12851 15351
rect 12851 15317 12860 15351
rect 12808 15308 12860 15317
rect 13176 15351 13228 15360
rect 13176 15317 13185 15351
rect 13185 15317 13219 15351
rect 13219 15317 13228 15351
rect 13176 15308 13228 15317
rect 13268 15351 13320 15360
rect 13268 15317 13277 15351
rect 13277 15317 13311 15351
rect 13311 15317 13320 15351
rect 13268 15308 13320 15317
rect 7898 15206 7950 15258
rect 7962 15206 8014 15258
rect 8026 15206 8078 15258
rect 8090 15206 8142 15258
rect 8154 15206 8206 15258
rect 14846 15206 14898 15258
rect 14910 15206 14962 15258
rect 14974 15206 15026 15258
rect 15038 15206 15090 15258
rect 15102 15206 15154 15258
rect 21794 15206 21846 15258
rect 21858 15206 21910 15258
rect 21922 15206 21974 15258
rect 21986 15206 22038 15258
rect 22050 15206 22102 15258
rect 4896 15147 4948 15156
rect 4896 15113 4905 15147
rect 4905 15113 4939 15147
rect 4939 15113 4948 15147
rect 4896 15104 4948 15113
rect 5448 15104 5500 15156
rect 13176 15104 13228 15156
rect 1952 14968 2004 15020
rect 2412 14968 2464 15020
rect 4160 14968 4212 15020
rect 6552 15011 6604 15020
rect 3608 14900 3660 14952
rect 6552 14977 6561 15011
rect 6561 14977 6595 15011
rect 6595 14977 6604 15011
rect 6552 14968 6604 14977
rect 11704 14968 11756 15020
rect 12164 14943 12216 14952
rect 12164 14909 12173 14943
rect 12173 14909 12207 14943
rect 12207 14909 12216 14943
rect 12164 14900 12216 14909
rect 2044 14764 2096 14816
rect 7748 14807 7800 14816
rect 7748 14773 7757 14807
rect 7757 14773 7791 14807
rect 7791 14773 7800 14807
rect 7748 14764 7800 14773
rect 27988 14764 28040 14816
rect 4424 14662 4476 14714
rect 4488 14662 4540 14714
rect 4552 14662 4604 14714
rect 4616 14662 4668 14714
rect 4680 14662 4732 14714
rect 11372 14662 11424 14714
rect 11436 14662 11488 14714
rect 11500 14662 11552 14714
rect 11564 14662 11616 14714
rect 11628 14662 11680 14714
rect 18320 14662 18372 14714
rect 18384 14662 18436 14714
rect 18448 14662 18500 14714
rect 18512 14662 18564 14714
rect 18576 14662 18628 14714
rect 25268 14662 25320 14714
rect 25332 14662 25384 14714
rect 25396 14662 25448 14714
rect 25460 14662 25512 14714
rect 25524 14662 25576 14714
rect 2872 14492 2924 14544
rect 3792 14492 3844 14544
rect 6552 14424 6604 14476
rect 9036 14560 9088 14612
rect 11796 14603 11848 14612
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3240 14356 3292 14365
rect 3792 14399 3844 14408
rect 3792 14365 3801 14399
rect 3801 14365 3835 14399
rect 3835 14365 3844 14399
rect 3792 14356 3844 14365
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 5080 14356 5132 14408
rect 7196 14356 7248 14408
rect 7288 14399 7340 14408
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7564 14399 7616 14408
rect 7288 14356 7340 14365
rect 7564 14365 7573 14399
rect 7573 14365 7607 14399
rect 7607 14365 7616 14399
rect 7564 14356 7616 14365
rect 10876 14492 10928 14544
rect 11796 14569 11805 14603
rect 11805 14569 11839 14603
rect 11839 14569 11848 14603
rect 11796 14560 11848 14569
rect 9496 14356 9548 14408
rect 10876 14356 10928 14408
rect 13268 14492 13320 14544
rect 11520 14467 11572 14476
rect 11520 14433 11529 14467
rect 11529 14433 11563 14467
rect 11563 14433 11572 14467
rect 11520 14424 11572 14433
rect 11428 14399 11480 14408
rect 11428 14365 11437 14399
rect 11437 14365 11471 14399
rect 11471 14365 11480 14399
rect 11428 14356 11480 14365
rect 2688 14288 2740 14340
rect 9864 14331 9916 14340
rect 9864 14297 9873 14331
rect 9873 14297 9907 14331
rect 9907 14297 9916 14331
rect 9864 14288 9916 14297
rect 11060 14288 11112 14340
rect 12532 14356 12584 14408
rect 12348 14331 12400 14340
rect 12348 14297 12357 14331
rect 12357 14297 12391 14331
rect 12391 14297 12400 14331
rect 12348 14288 12400 14297
rect 2136 14263 2188 14272
rect 2136 14229 2145 14263
rect 2145 14229 2179 14263
rect 2179 14229 2188 14263
rect 2136 14220 2188 14229
rect 2780 14220 2832 14272
rect 3884 14263 3936 14272
rect 3884 14229 3893 14263
rect 3893 14229 3927 14263
rect 3927 14229 3936 14263
rect 3884 14220 3936 14229
rect 3976 14220 4028 14272
rect 6460 14263 6512 14272
rect 6460 14229 6469 14263
rect 6469 14229 6503 14263
rect 6503 14229 6512 14263
rect 6460 14220 6512 14229
rect 7288 14220 7340 14272
rect 9680 14220 9732 14272
rect 10048 14220 10100 14272
rect 12256 14220 12308 14272
rect 7898 14118 7950 14170
rect 7962 14118 8014 14170
rect 8026 14118 8078 14170
rect 8090 14118 8142 14170
rect 8154 14118 8206 14170
rect 14846 14118 14898 14170
rect 14910 14118 14962 14170
rect 14974 14118 15026 14170
rect 15038 14118 15090 14170
rect 15102 14118 15154 14170
rect 21794 14118 21846 14170
rect 21858 14118 21910 14170
rect 21922 14118 21974 14170
rect 21986 14118 22038 14170
rect 22050 14118 22102 14170
rect 3240 14016 3292 14068
rect 7748 14016 7800 14068
rect 8760 14059 8812 14068
rect 8760 14025 8769 14059
rect 8769 14025 8803 14059
rect 8803 14025 8812 14059
rect 8760 14016 8812 14025
rect 9588 14016 9640 14068
rect 12992 14059 13044 14068
rect 12992 14025 13001 14059
rect 13001 14025 13035 14059
rect 13035 14025 13044 14059
rect 12992 14016 13044 14025
rect 1676 13855 1728 13864
rect 1676 13821 1685 13855
rect 1685 13821 1719 13855
rect 1719 13821 1728 13855
rect 1676 13812 1728 13821
rect 2872 13923 2924 13932
rect 2872 13889 2881 13923
rect 2881 13889 2915 13923
rect 2915 13889 2924 13923
rect 3148 13948 3200 14000
rect 4068 13948 4120 14000
rect 2872 13880 2924 13889
rect 3884 13923 3936 13932
rect 3884 13889 3893 13923
rect 3893 13889 3927 13923
rect 3927 13889 3936 13923
rect 3884 13880 3936 13889
rect 6644 13948 6696 14000
rect 9680 13948 9732 14000
rect 11428 13948 11480 14000
rect 6552 13880 6604 13932
rect 3240 13812 3292 13864
rect 3608 13855 3660 13864
rect 3608 13821 3617 13855
rect 3617 13821 3651 13855
rect 3651 13821 3660 13855
rect 3608 13812 3660 13821
rect 6736 13812 6788 13864
rect 9128 13880 9180 13932
rect 9772 13880 9824 13932
rect 12348 13880 12400 13932
rect 13728 13880 13780 13932
rect 1952 13787 2004 13796
rect 1952 13753 1961 13787
rect 1961 13753 1995 13787
rect 1995 13753 2004 13787
rect 1952 13744 2004 13753
rect 2964 13787 3016 13796
rect 2964 13753 2973 13787
rect 2973 13753 3007 13787
rect 3007 13753 3016 13787
rect 2964 13744 3016 13753
rect 5816 13787 5868 13796
rect 5816 13753 5825 13787
rect 5825 13753 5859 13787
rect 5859 13753 5868 13787
rect 5816 13744 5868 13753
rect 6828 13744 6880 13796
rect 9312 13812 9364 13864
rect 9864 13812 9916 13864
rect 9956 13855 10008 13864
rect 9956 13821 9965 13855
rect 9965 13821 9999 13855
rect 9999 13821 10008 13855
rect 9956 13812 10008 13821
rect 11520 13812 11572 13864
rect 13820 13812 13872 13864
rect 7472 13676 7524 13728
rect 9404 13744 9456 13796
rect 11888 13744 11940 13796
rect 14096 13744 14148 13796
rect 10048 13676 10100 13728
rect 11060 13676 11112 13728
rect 13268 13719 13320 13728
rect 13268 13685 13277 13719
rect 13277 13685 13311 13719
rect 13311 13685 13320 13719
rect 13268 13676 13320 13685
rect 4424 13574 4476 13626
rect 4488 13574 4540 13626
rect 4552 13574 4604 13626
rect 4616 13574 4668 13626
rect 4680 13574 4732 13626
rect 11372 13574 11424 13626
rect 11436 13574 11488 13626
rect 11500 13574 11552 13626
rect 11564 13574 11616 13626
rect 11628 13574 11680 13626
rect 18320 13574 18372 13626
rect 18384 13574 18436 13626
rect 18448 13574 18500 13626
rect 18512 13574 18564 13626
rect 18576 13574 18628 13626
rect 25268 13574 25320 13626
rect 25332 13574 25384 13626
rect 25396 13574 25448 13626
rect 25460 13574 25512 13626
rect 25524 13574 25576 13626
rect 1952 13472 2004 13524
rect 9772 13472 9824 13524
rect 9956 13404 10008 13456
rect 13820 13472 13872 13524
rect 15568 13472 15620 13524
rect 10876 13404 10928 13456
rect 2688 13379 2740 13388
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 2688 13345 2697 13379
rect 2697 13345 2731 13379
rect 2731 13345 2740 13379
rect 2688 13336 2740 13345
rect 3148 13336 3200 13388
rect 6368 13336 6420 13388
rect 6828 13379 6880 13388
rect 6828 13345 6837 13379
rect 6837 13345 6871 13379
rect 6871 13345 6880 13379
rect 6828 13336 6880 13345
rect 5080 13311 5132 13320
rect 1768 13175 1820 13184
rect 1768 13141 1777 13175
rect 1777 13141 1811 13175
rect 1811 13141 1820 13175
rect 1768 13132 1820 13141
rect 5080 13277 5089 13311
rect 5089 13277 5123 13311
rect 5123 13277 5132 13311
rect 5080 13268 5132 13277
rect 9772 13336 9824 13388
rect 11060 13336 11112 13388
rect 12348 13336 12400 13388
rect 2872 13200 2924 13252
rect 4252 13243 4304 13252
rect 4252 13209 4261 13243
rect 4261 13209 4295 13243
rect 4295 13209 4304 13243
rect 4252 13200 4304 13209
rect 9404 13268 9456 13320
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 11244 13268 11296 13320
rect 12808 13268 12860 13320
rect 14372 13311 14424 13320
rect 14372 13277 14381 13311
rect 14381 13277 14415 13311
rect 14415 13277 14424 13311
rect 14372 13268 14424 13277
rect 9864 13243 9916 13252
rect 9864 13209 9873 13243
rect 9873 13209 9907 13243
rect 9907 13209 9916 13243
rect 9864 13200 9916 13209
rect 14188 13200 14240 13252
rect 15292 13268 15344 13320
rect 2964 13132 3016 13184
rect 4988 13175 5040 13184
rect 4988 13141 4997 13175
rect 4997 13141 5031 13175
rect 5031 13141 5040 13175
rect 4988 13132 5040 13141
rect 5448 13132 5500 13184
rect 6184 13175 6236 13184
rect 6184 13141 6193 13175
rect 6193 13141 6227 13175
rect 6227 13141 6236 13175
rect 6184 13132 6236 13141
rect 6552 13175 6604 13184
rect 6552 13141 6561 13175
rect 6561 13141 6595 13175
rect 6595 13141 6604 13175
rect 6552 13132 6604 13141
rect 7656 13132 7708 13184
rect 10692 13132 10744 13184
rect 10784 13132 10836 13184
rect 11980 13175 12032 13184
rect 11980 13141 11989 13175
rect 11989 13141 12023 13175
rect 12023 13141 12032 13175
rect 11980 13132 12032 13141
rect 12532 13132 12584 13184
rect 7898 13030 7950 13082
rect 7962 13030 8014 13082
rect 8026 13030 8078 13082
rect 8090 13030 8142 13082
rect 8154 13030 8206 13082
rect 14846 13030 14898 13082
rect 14910 13030 14962 13082
rect 14974 13030 15026 13082
rect 15038 13030 15090 13082
rect 15102 13030 15154 13082
rect 21794 13030 21846 13082
rect 21858 13030 21910 13082
rect 21922 13030 21974 13082
rect 21986 13030 22038 13082
rect 22050 13030 22102 13082
rect 2688 12928 2740 12980
rect 4252 12928 4304 12980
rect 14372 12928 14424 12980
rect 2872 12860 2924 12912
rect 2964 12792 3016 12844
rect 3332 12792 3384 12844
rect 5080 12792 5132 12844
rect 7472 12835 7524 12844
rect 3516 12724 3568 12776
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 9772 12792 9824 12844
rect 10876 12792 10928 12844
rect 11980 12835 12032 12844
rect 11980 12801 11989 12835
rect 11989 12801 12023 12835
rect 12023 12801 12032 12835
rect 11980 12792 12032 12801
rect 14188 12792 14240 12844
rect 13636 12724 13688 12776
rect 2412 12699 2464 12708
rect 2412 12665 2421 12699
rect 2421 12665 2455 12699
rect 2455 12665 2464 12699
rect 2412 12656 2464 12665
rect 3884 12656 3936 12708
rect 15568 12656 15620 12708
rect 4804 12588 4856 12640
rect 6920 12631 6972 12640
rect 6920 12597 6929 12631
rect 6929 12597 6963 12631
rect 6963 12597 6972 12631
rect 6920 12588 6972 12597
rect 7748 12588 7800 12640
rect 9680 12588 9732 12640
rect 11796 12631 11848 12640
rect 11796 12597 11805 12631
rect 11805 12597 11839 12631
rect 11839 12597 11848 12631
rect 11796 12588 11848 12597
rect 13912 12631 13964 12640
rect 13912 12597 13921 12631
rect 13921 12597 13955 12631
rect 13955 12597 13964 12631
rect 13912 12588 13964 12597
rect 4424 12486 4476 12538
rect 4488 12486 4540 12538
rect 4552 12486 4604 12538
rect 4616 12486 4668 12538
rect 4680 12486 4732 12538
rect 11372 12486 11424 12538
rect 11436 12486 11488 12538
rect 11500 12486 11552 12538
rect 11564 12486 11616 12538
rect 11628 12486 11680 12538
rect 18320 12486 18372 12538
rect 18384 12486 18436 12538
rect 18448 12486 18500 12538
rect 18512 12486 18564 12538
rect 18576 12486 18628 12538
rect 25268 12486 25320 12538
rect 25332 12486 25384 12538
rect 25396 12486 25448 12538
rect 25460 12486 25512 12538
rect 25524 12486 25576 12538
rect 12348 12248 12400 12300
rect 6184 12180 6236 12232
rect 12532 12180 12584 12232
rect 13268 12180 13320 12232
rect 18144 12384 18196 12436
rect 4252 12044 4304 12096
rect 14740 12044 14792 12096
rect 7898 11942 7950 11994
rect 7962 11942 8014 11994
rect 8026 11942 8078 11994
rect 8090 11942 8142 11994
rect 8154 11942 8206 11994
rect 14846 11942 14898 11994
rect 14910 11942 14962 11994
rect 14974 11942 15026 11994
rect 15038 11942 15090 11994
rect 15102 11942 15154 11994
rect 21794 11942 21846 11994
rect 21858 11942 21910 11994
rect 21922 11942 21974 11994
rect 21986 11942 22038 11994
rect 22050 11942 22102 11994
rect 9864 11840 9916 11892
rect 14832 11704 14884 11756
rect 4344 11500 4396 11552
rect 11796 11636 11848 11688
rect 8484 11500 8536 11552
rect 10600 11500 10652 11552
rect 11704 11543 11756 11552
rect 11704 11509 11713 11543
rect 11713 11509 11747 11543
rect 11747 11509 11756 11543
rect 11704 11500 11756 11509
rect 4424 11398 4476 11450
rect 4488 11398 4540 11450
rect 4552 11398 4604 11450
rect 4616 11398 4668 11450
rect 4680 11398 4732 11450
rect 11372 11398 11424 11450
rect 11436 11398 11488 11450
rect 11500 11398 11552 11450
rect 11564 11398 11616 11450
rect 11628 11398 11680 11450
rect 18320 11398 18372 11450
rect 18384 11398 18436 11450
rect 18448 11398 18500 11450
rect 18512 11398 18564 11450
rect 18576 11398 18628 11450
rect 25268 11398 25320 11450
rect 25332 11398 25384 11450
rect 25396 11398 25448 11450
rect 25460 11398 25512 11450
rect 25524 11398 25576 11450
rect 3148 11296 3200 11348
rect 6368 11296 6420 11348
rect 13636 11296 13688 11348
rect 14832 11339 14884 11348
rect 14832 11305 14841 11339
rect 14841 11305 14875 11339
rect 14875 11305 14884 11339
rect 14832 11296 14884 11305
rect 2780 11160 2832 11212
rect 1492 11135 1544 11144
rect 1492 11101 1501 11135
rect 1501 11101 1535 11135
rect 1535 11101 1544 11135
rect 1492 11092 1544 11101
rect 3976 11228 4028 11280
rect 4252 11203 4304 11212
rect 4252 11169 4261 11203
rect 4261 11169 4295 11203
rect 4295 11169 4304 11203
rect 4252 11160 4304 11169
rect 13912 11160 13964 11212
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 10324 11092 10376 11144
rect 14096 11092 14148 11144
rect 14648 11092 14700 11144
rect 4804 11024 4856 11076
rect 9680 11024 9732 11076
rect 7898 10854 7950 10906
rect 7962 10854 8014 10906
rect 8026 10854 8078 10906
rect 8090 10854 8142 10906
rect 8154 10854 8206 10906
rect 14846 10854 14898 10906
rect 14910 10854 14962 10906
rect 14974 10854 15026 10906
rect 15038 10854 15090 10906
rect 15102 10854 15154 10906
rect 21794 10854 21846 10906
rect 21858 10854 21910 10906
rect 21922 10854 21974 10906
rect 21986 10854 22038 10906
rect 22050 10854 22102 10906
rect 1492 10752 1544 10804
rect 3976 10752 4028 10804
rect 9036 10795 9088 10804
rect 9036 10761 9045 10795
rect 9045 10761 9079 10795
rect 9079 10761 9088 10795
rect 9036 10752 9088 10761
rect 13268 10795 13320 10804
rect 13268 10761 13277 10795
rect 13277 10761 13311 10795
rect 13311 10761 13320 10795
rect 13268 10752 13320 10761
rect 2136 10727 2188 10736
rect 2136 10693 2145 10727
rect 2145 10693 2179 10727
rect 2179 10693 2188 10727
rect 2136 10684 2188 10693
rect 3884 10684 3936 10736
rect 4344 10727 4396 10736
rect 4344 10693 4353 10727
rect 4353 10693 4387 10727
rect 4387 10693 4396 10727
rect 4344 10684 4396 10693
rect 7288 10684 7340 10736
rect 9496 10684 9548 10736
rect 10784 10684 10836 10736
rect 13728 10684 13780 10736
rect 5448 10616 5500 10668
rect 5816 10616 5868 10668
rect 14740 10616 14792 10668
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 6368 10591 6420 10600
rect 6368 10557 6377 10591
rect 6377 10557 6411 10591
rect 6411 10557 6420 10591
rect 6368 10548 6420 10557
rect 6644 10548 6696 10600
rect 4160 10412 4212 10464
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 5816 10412 5868 10421
rect 10324 10412 10376 10464
rect 4424 10310 4476 10362
rect 4488 10310 4540 10362
rect 4552 10310 4604 10362
rect 4616 10310 4668 10362
rect 4680 10310 4732 10362
rect 11372 10310 11424 10362
rect 11436 10310 11488 10362
rect 11500 10310 11552 10362
rect 11564 10310 11616 10362
rect 11628 10310 11680 10362
rect 18320 10310 18372 10362
rect 18384 10310 18436 10362
rect 18448 10310 18500 10362
rect 18512 10310 18564 10362
rect 18576 10310 18628 10362
rect 25268 10310 25320 10362
rect 25332 10310 25384 10362
rect 25396 10310 25448 10362
rect 25460 10310 25512 10362
rect 25524 10310 25576 10362
rect 3240 10251 3292 10260
rect 3240 10217 3249 10251
rect 3249 10217 3283 10251
rect 3283 10217 3292 10251
rect 3240 10208 3292 10217
rect 5816 10208 5868 10260
rect 14004 10208 14056 10260
rect 7380 10140 7432 10192
rect 1768 10115 1820 10124
rect 1768 10081 1777 10115
rect 1777 10081 1811 10115
rect 1811 10081 1820 10115
rect 1768 10072 1820 10081
rect 6368 10072 6420 10124
rect 6460 10072 6512 10124
rect 10600 10115 10652 10124
rect 10600 10081 10609 10115
rect 10609 10081 10643 10115
rect 10643 10081 10652 10115
rect 10600 10072 10652 10081
rect 11152 10072 11204 10124
rect 1492 10047 1544 10056
rect 1492 10013 1501 10047
rect 1501 10013 1535 10047
rect 1535 10013 1544 10047
rect 1492 10004 1544 10013
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 14648 10047 14700 10056
rect 14648 10013 14657 10047
rect 14657 10013 14691 10047
rect 14691 10013 14700 10047
rect 14648 10004 14700 10013
rect 3516 9936 3568 9988
rect 6920 9936 6972 9988
rect 12716 9936 12768 9988
rect 13728 9868 13780 9920
rect 7898 9766 7950 9818
rect 7962 9766 8014 9818
rect 8026 9766 8078 9818
rect 8090 9766 8142 9818
rect 8154 9766 8206 9818
rect 14846 9766 14898 9818
rect 14910 9766 14962 9818
rect 14974 9766 15026 9818
rect 15038 9766 15090 9818
rect 15102 9766 15154 9818
rect 21794 9766 21846 9818
rect 21858 9766 21910 9818
rect 21922 9766 21974 9818
rect 21986 9766 22038 9818
rect 22050 9766 22102 9818
rect 2044 9639 2096 9648
rect 2044 9605 2053 9639
rect 2053 9605 2087 9639
rect 2087 9605 2096 9639
rect 2044 9596 2096 9605
rect 4988 9596 5040 9648
rect 11152 9596 11204 9648
rect 11704 9596 11756 9648
rect 13728 9596 13780 9648
rect 8484 9528 8536 9580
rect 10324 9528 10376 9580
rect 14648 9596 14700 9648
rect 1492 9460 1544 9512
rect 3332 9460 3384 9512
rect 6552 9460 6604 9512
rect 7748 9460 7800 9512
rect 10692 9460 10744 9512
rect 15292 9571 15344 9580
rect 15292 9537 15301 9571
rect 15301 9537 15335 9571
rect 15335 9537 15344 9571
rect 15292 9528 15344 9537
rect 14280 9460 14332 9512
rect 3240 9324 3292 9376
rect 14004 9367 14056 9376
rect 14004 9333 14013 9367
rect 14013 9333 14047 9367
rect 14047 9333 14056 9367
rect 14004 9324 14056 9333
rect 15384 9324 15436 9376
rect 16672 9367 16724 9376
rect 16672 9333 16681 9367
rect 16681 9333 16715 9367
rect 16715 9333 16724 9367
rect 16672 9324 16724 9333
rect 18972 9367 19024 9376
rect 18972 9333 18981 9367
rect 18981 9333 19015 9367
rect 19015 9333 19024 9367
rect 18972 9324 19024 9333
rect 19616 9367 19668 9376
rect 19616 9333 19625 9367
rect 19625 9333 19659 9367
rect 19659 9333 19668 9367
rect 19616 9324 19668 9333
rect 4424 9222 4476 9274
rect 4488 9222 4540 9274
rect 4552 9222 4604 9274
rect 4616 9222 4668 9274
rect 4680 9222 4732 9274
rect 11372 9222 11424 9274
rect 11436 9222 11488 9274
rect 11500 9222 11552 9274
rect 11564 9222 11616 9274
rect 11628 9222 11680 9274
rect 18320 9222 18372 9274
rect 18384 9222 18436 9274
rect 18448 9222 18500 9274
rect 18512 9222 18564 9274
rect 18576 9222 18628 9274
rect 25268 9222 25320 9274
rect 25332 9222 25384 9274
rect 25396 9222 25448 9274
rect 25460 9222 25512 9274
rect 25524 9222 25576 9274
rect 7564 9120 7616 9172
rect 12716 9120 12768 9172
rect 3240 8984 3292 9036
rect 4068 8984 4120 9036
rect 6368 8984 6420 9036
rect 6644 8984 6696 9036
rect 7012 8984 7064 9036
rect 7564 8984 7616 9036
rect 19616 9120 19668 9172
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 14740 8916 14792 8968
rect 6552 8848 6604 8900
rect 7656 8848 7708 8900
rect 7898 8678 7950 8730
rect 7962 8678 8014 8730
rect 8026 8678 8078 8730
rect 8090 8678 8142 8730
rect 8154 8678 8206 8730
rect 14846 8678 14898 8730
rect 14910 8678 14962 8730
rect 14974 8678 15026 8730
rect 15038 8678 15090 8730
rect 15102 8678 15154 8730
rect 21794 8678 21846 8730
rect 21858 8678 21910 8730
rect 21922 8678 21974 8730
rect 21986 8678 22038 8730
rect 22050 8678 22102 8730
rect 4804 8508 4856 8560
rect 9772 8508 9824 8560
rect 12348 8508 12400 8560
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 8484 8440 8536 8492
rect 14740 8440 14792 8492
rect 3516 8415 3568 8424
rect 3516 8381 3525 8415
rect 3525 8381 3559 8415
rect 3559 8381 3568 8415
rect 3516 8372 3568 8381
rect 14004 8415 14056 8424
rect 14004 8381 14013 8415
rect 14013 8381 14047 8415
rect 14047 8381 14056 8415
rect 14004 8372 14056 8381
rect 6276 8304 6328 8356
rect 6644 8304 6696 8356
rect 14096 8304 14148 8356
rect 11244 8236 11296 8288
rect 4424 8134 4476 8186
rect 4488 8134 4540 8186
rect 4552 8134 4604 8186
rect 4616 8134 4668 8186
rect 4680 8134 4732 8186
rect 11372 8134 11424 8186
rect 11436 8134 11488 8186
rect 11500 8134 11552 8186
rect 11564 8134 11616 8186
rect 11628 8134 11680 8186
rect 18320 8134 18372 8186
rect 18384 8134 18436 8186
rect 18448 8134 18500 8186
rect 18512 8134 18564 8186
rect 18576 8134 18628 8186
rect 25268 8134 25320 8186
rect 25332 8134 25384 8186
rect 25396 8134 25448 8186
rect 25460 8134 25512 8186
rect 25524 8134 25576 8186
rect 3516 8032 3568 8084
rect 9772 8075 9824 8084
rect 9772 8041 9781 8075
rect 9781 8041 9815 8075
rect 9815 8041 9824 8075
rect 9772 8032 9824 8041
rect 12348 8032 12400 8084
rect 14096 8075 14148 8084
rect 14096 8041 14105 8075
rect 14105 8041 14139 8075
rect 14139 8041 14148 8075
rect 14096 8032 14148 8041
rect 15568 8075 15620 8084
rect 15568 8041 15577 8075
rect 15577 8041 15611 8075
rect 15611 8041 15620 8075
rect 15568 8032 15620 8041
rect 3240 7896 3292 7948
rect 8484 7896 8536 7948
rect 11244 7896 11296 7948
rect 11336 7896 11388 7948
rect 1768 7803 1820 7812
rect 1768 7769 1777 7803
rect 1777 7769 1811 7803
rect 1811 7769 1820 7803
rect 1768 7760 1820 7769
rect 3700 7760 3752 7812
rect 4344 7760 4396 7812
rect 7656 7760 7708 7812
rect 12256 7760 12308 7812
rect 4896 7692 4948 7744
rect 6184 7735 6236 7744
rect 6184 7701 6193 7735
rect 6193 7701 6227 7735
rect 6227 7701 6236 7735
rect 6184 7692 6236 7701
rect 14280 7828 14332 7880
rect 14464 7828 14516 7880
rect 15384 7871 15436 7880
rect 15384 7837 15393 7871
rect 15393 7837 15427 7871
rect 15427 7837 15436 7871
rect 15384 7828 15436 7837
rect 14740 7760 14792 7812
rect 16672 7803 16724 7812
rect 16672 7769 16681 7803
rect 16681 7769 16715 7803
rect 16715 7769 16724 7803
rect 16672 7760 16724 7769
rect 23296 7692 23348 7744
rect 7898 7590 7950 7642
rect 7962 7590 8014 7642
rect 8026 7590 8078 7642
rect 8090 7590 8142 7642
rect 8154 7590 8206 7642
rect 14846 7590 14898 7642
rect 14910 7590 14962 7642
rect 14974 7590 15026 7642
rect 15038 7590 15090 7642
rect 15102 7590 15154 7642
rect 21794 7590 21846 7642
rect 21858 7590 21910 7642
rect 21922 7590 21974 7642
rect 21986 7590 22038 7642
rect 22050 7590 22102 7642
rect 3240 7488 3292 7540
rect 11336 7488 11388 7540
rect 12256 7488 12308 7540
rect 6184 7420 6236 7472
rect 14004 7420 14056 7472
rect 1768 7352 1820 7404
rect 4344 7395 4396 7404
rect 4344 7361 4353 7395
rect 4353 7361 4387 7395
rect 4387 7361 4396 7395
rect 4344 7352 4396 7361
rect 8484 7352 8536 7404
rect 10048 7284 10100 7336
rect 14740 7352 14792 7404
rect 14648 7284 14700 7336
rect 10784 7216 10836 7268
rect 4988 7191 5040 7200
rect 4988 7157 4997 7191
rect 4997 7157 5031 7191
rect 5031 7157 5040 7191
rect 4988 7148 5040 7157
rect 5816 7191 5868 7200
rect 5816 7157 5825 7191
rect 5825 7157 5859 7191
rect 5859 7157 5868 7191
rect 5816 7148 5868 7157
rect 7656 7148 7708 7200
rect 13176 7148 13228 7200
rect 4424 7046 4476 7098
rect 4488 7046 4540 7098
rect 4552 7046 4604 7098
rect 4616 7046 4668 7098
rect 4680 7046 4732 7098
rect 11372 7046 11424 7098
rect 11436 7046 11488 7098
rect 11500 7046 11552 7098
rect 11564 7046 11616 7098
rect 11628 7046 11680 7098
rect 18320 7046 18372 7098
rect 18384 7046 18436 7098
rect 18448 7046 18500 7098
rect 18512 7046 18564 7098
rect 18576 7046 18628 7098
rect 25268 7046 25320 7098
rect 25332 7046 25384 7098
rect 25396 7046 25448 7098
rect 25460 7046 25512 7098
rect 25524 7046 25576 7098
rect 4988 6944 5040 6996
rect 5816 6944 5868 6996
rect 14096 6987 14148 6996
rect 14096 6953 14105 6987
rect 14105 6953 14139 6987
rect 14139 6953 14148 6987
rect 14096 6944 14148 6953
rect 6736 6808 6788 6860
rect 10784 6808 10836 6860
rect 11244 6808 11296 6860
rect 2320 6783 2372 6792
rect 2320 6749 2329 6783
rect 2329 6749 2363 6783
rect 2363 6749 2372 6783
rect 2320 6740 2372 6749
rect 3148 6783 3200 6792
rect 3148 6749 3157 6783
rect 3157 6749 3191 6783
rect 3191 6749 3200 6783
rect 3148 6740 3200 6749
rect 3608 6740 3660 6792
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 10324 6740 10376 6792
rect 14372 6783 14424 6792
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 15200 6740 15252 6792
rect 6736 6672 6788 6724
rect 10692 6672 10744 6724
rect 11152 6715 11204 6724
rect 11152 6681 11161 6715
rect 11161 6681 11195 6715
rect 11195 6681 11204 6715
rect 11152 6672 11204 6681
rect 13176 6672 13228 6724
rect 14096 6715 14148 6724
rect 14096 6681 14105 6715
rect 14105 6681 14139 6715
rect 14139 6681 14148 6715
rect 14096 6672 14148 6681
rect 3056 6647 3108 6656
rect 3056 6613 3065 6647
rect 3065 6613 3099 6647
rect 3099 6613 3108 6647
rect 3056 6604 3108 6613
rect 5908 6647 5960 6656
rect 5908 6613 5917 6647
rect 5917 6613 5951 6647
rect 5951 6613 5960 6647
rect 5908 6604 5960 6613
rect 6552 6604 6604 6656
rect 12808 6604 12860 6656
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 16580 6647 16632 6656
rect 16580 6613 16589 6647
rect 16589 6613 16623 6647
rect 16623 6613 16632 6647
rect 16580 6604 16632 6613
rect 7898 6502 7950 6554
rect 7962 6502 8014 6554
rect 8026 6502 8078 6554
rect 8090 6502 8142 6554
rect 8154 6502 8206 6554
rect 14846 6502 14898 6554
rect 14910 6502 14962 6554
rect 14974 6502 15026 6554
rect 15038 6502 15090 6554
rect 15102 6502 15154 6554
rect 21794 6502 21846 6554
rect 21858 6502 21910 6554
rect 21922 6502 21974 6554
rect 21986 6502 22038 6554
rect 22050 6502 22102 6554
rect 4804 6400 4856 6452
rect 11244 6400 11296 6452
rect 14188 6443 14240 6452
rect 2320 6375 2372 6384
rect 2320 6341 2329 6375
rect 2329 6341 2363 6375
rect 2363 6341 2372 6375
rect 2320 6332 2372 6341
rect 3608 6332 3660 6384
rect 5356 6375 5408 6384
rect 3424 6264 3476 6316
rect 5356 6341 5365 6375
rect 5365 6341 5399 6375
rect 5399 6341 5408 6375
rect 5356 6332 5408 6341
rect 6644 6375 6696 6384
rect 6644 6341 6653 6375
rect 6653 6341 6687 6375
rect 6687 6341 6696 6375
rect 6644 6332 6696 6341
rect 12808 6375 12860 6384
rect 12808 6341 12817 6375
rect 12817 6341 12851 6375
rect 12851 6341 12860 6375
rect 12808 6332 12860 6341
rect 14188 6409 14197 6443
rect 14197 6409 14231 6443
rect 14231 6409 14240 6443
rect 14188 6400 14240 6409
rect 14648 6400 14700 6452
rect 14464 6332 14516 6384
rect 7748 6264 7800 6316
rect 11060 6264 11112 6316
rect 11152 6264 11204 6316
rect 8576 6239 8628 6248
rect 8576 6205 8585 6239
rect 8585 6205 8619 6239
rect 8619 6205 8628 6239
rect 8576 6196 8628 6205
rect 8944 6196 8996 6248
rect 13176 6264 13228 6316
rect 14004 6307 14056 6316
rect 14004 6273 14013 6307
rect 14013 6273 14047 6307
rect 14047 6273 14056 6307
rect 14004 6264 14056 6273
rect 15200 6264 15252 6316
rect 12900 6239 12952 6248
rect 12900 6205 12909 6239
rect 12909 6205 12943 6239
rect 12943 6205 12952 6239
rect 12900 6196 12952 6205
rect 2780 6060 2832 6112
rect 3792 6103 3844 6112
rect 3792 6069 3801 6103
rect 3801 6069 3835 6103
rect 3835 6069 3844 6103
rect 3792 6060 3844 6069
rect 8668 6060 8720 6112
rect 12808 6103 12860 6112
rect 12808 6069 12817 6103
rect 12817 6069 12851 6103
rect 12851 6069 12860 6103
rect 12808 6060 12860 6069
rect 14556 6060 14608 6112
rect 4424 5958 4476 6010
rect 4488 5958 4540 6010
rect 4552 5958 4604 6010
rect 4616 5958 4668 6010
rect 4680 5958 4732 6010
rect 11372 5958 11424 6010
rect 11436 5958 11488 6010
rect 11500 5958 11552 6010
rect 11564 5958 11616 6010
rect 11628 5958 11680 6010
rect 18320 5958 18372 6010
rect 18384 5958 18436 6010
rect 18448 5958 18500 6010
rect 18512 5958 18564 6010
rect 18576 5958 18628 6010
rect 25268 5958 25320 6010
rect 25332 5958 25384 6010
rect 25396 5958 25448 6010
rect 25460 5958 25512 6010
rect 25524 5958 25576 6010
rect 3792 5856 3844 5908
rect 8668 5856 8720 5908
rect 8944 5899 8996 5908
rect 8944 5865 8953 5899
rect 8953 5865 8987 5899
rect 8987 5865 8996 5899
rect 8944 5856 8996 5865
rect 12808 5856 12860 5908
rect 11060 5788 11112 5840
rect 6552 5763 6604 5772
rect 6552 5729 6561 5763
rect 6561 5729 6595 5763
rect 6595 5729 6604 5763
rect 6552 5720 6604 5729
rect 8576 5720 8628 5772
rect 10324 5720 10376 5772
rect 10692 5720 10744 5772
rect 6276 5652 6328 5704
rect 7472 5652 7524 5704
rect 9956 5627 10008 5636
rect 9956 5593 9965 5627
rect 9965 5593 9999 5627
rect 9999 5593 10008 5627
rect 9956 5584 10008 5593
rect 13084 5584 13136 5636
rect 15200 5652 15252 5704
rect 13544 5516 13596 5568
rect 14740 5516 14792 5568
rect 7898 5414 7950 5466
rect 7962 5414 8014 5466
rect 8026 5414 8078 5466
rect 8090 5414 8142 5466
rect 8154 5414 8206 5466
rect 14846 5414 14898 5466
rect 14910 5414 14962 5466
rect 14974 5414 15026 5466
rect 15038 5414 15090 5466
rect 15102 5414 15154 5466
rect 21794 5414 21846 5466
rect 21858 5414 21910 5466
rect 21922 5414 21974 5466
rect 21986 5414 22038 5466
rect 22050 5414 22102 5466
rect 8576 5312 8628 5364
rect 5264 5219 5316 5228
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 3792 5108 3844 5160
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 7656 5244 7708 5296
rect 19892 5244 19944 5296
rect 9956 5176 10008 5228
rect 14280 5176 14332 5228
rect 14648 5176 14700 5228
rect 5080 5151 5132 5160
rect 5080 5117 5089 5151
rect 5089 5117 5123 5151
rect 5123 5117 5132 5151
rect 5080 5108 5132 5117
rect 8116 5108 8168 5160
rect 14096 5108 14148 5160
rect 13176 5040 13228 5092
rect 1768 4972 1820 5024
rect 4896 4972 4948 5024
rect 6644 4972 6696 5024
rect 11704 5015 11756 5024
rect 11704 4981 11713 5015
rect 11713 4981 11747 5015
rect 11747 4981 11756 5015
rect 11704 4972 11756 4981
rect 13728 5015 13780 5024
rect 13728 4981 13737 5015
rect 13737 4981 13771 5015
rect 13771 4981 13780 5015
rect 13728 4972 13780 4981
rect 4424 4870 4476 4922
rect 4488 4870 4540 4922
rect 4552 4870 4604 4922
rect 4616 4870 4668 4922
rect 4680 4870 4732 4922
rect 11372 4870 11424 4922
rect 11436 4870 11488 4922
rect 11500 4870 11552 4922
rect 11564 4870 11616 4922
rect 11628 4870 11680 4922
rect 18320 4870 18372 4922
rect 18384 4870 18436 4922
rect 18448 4870 18500 4922
rect 18512 4870 18564 4922
rect 18576 4870 18628 4922
rect 25268 4870 25320 4922
rect 25332 4870 25384 4922
rect 25396 4870 25448 4922
rect 25460 4870 25512 4922
rect 25524 4870 25576 4922
rect 3792 4811 3844 4820
rect 3792 4777 3801 4811
rect 3801 4777 3835 4811
rect 3835 4777 3844 4811
rect 3792 4768 3844 4777
rect 8116 4811 8168 4820
rect 8116 4777 8125 4811
rect 8125 4777 8159 4811
rect 8159 4777 8168 4811
rect 8116 4768 8168 4777
rect 13084 4768 13136 4820
rect 14188 4768 14240 4820
rect 16580 4768 16632 4820
rect 19892 4811 19944 4820
rect 19892 4777 19901 4811
rect 19901 4777 19935 4811
rect 19935 4777 19944 4811
rect 19892 4768 19944 4777
rect 5080 4700 5132 4752
rect 2780 4632 2832 4684
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 6644 4675 6696 4684
rect 6644 4641 6653 4675
rect 6653 4641 6687 4675
rect 6687 4641 6696 4675
rect 6644 4632 6696 4641
rect 10324 4675 10376 4684
rect 10324 4641 10333 4675
rect 10333 4641 10367 4675
rect 10367 4641 10376 4675
rect 10324 4632 10376 4641
rect 10968 4632 11020 4684
rect 4160 4564 4212 4616
rect 4896 4564 4948 4616
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 1768 4539 1820 4548
rect 1768 4505 1777 4539
rect 1777 4505 1811 4539
rect 1811 4505 1820 4539
rect 1768 4496 1820 4505
rect 3056 4496 3108 4548
rect 7656 4496 7708 4548
rect 10600 4539 10652 4548
rect 10600 4505 10609 4539
rect 10609 4505 10643 4539
rect 10643 4505 10652 4539
rect 10600 4496 10652 4505
rect 4620 4471 4672 4480
rect 4620 4437 4629 4471
rect 4629 4437 4663 4471
rect 4663 4437 4672 4471
rect 4620 4428 4672 4437
rect 13544 4428 13596 4480
rect 16580 4564 16632 4616
rect 16212 4496 16264 4548
rect 16396 4471 16448 4480
rect 16396 4437 16405 4471
rect 16405 4437 16439 4471
rect 16439 4437 16448 4471
rect 16396 4428 16448 4437
rect 7898 4326 7950 4378
rect 7962 4326 8014 4378
rect 8026 4326 8078 4378
rect 8090 4326 8142 4378
rect 8154 4326 8206 4378
rect 14846 4326 14898 4378
rect 14910 4326 14962 4378
rect 14974 4326 15026 4378
rect 15038 4326 15090 4378
rect 15102 4326 15154 4378
rect 21794 4326 21846 4378
rect 21858 4326 21910 4378
rect 21922 4326 21974 4378
rect 21986 4326 22038 4378
rect 22050 4326 22102 4378
rect 4620 4156 4672 4208
rect 16120 4224 16172 4276
rect 11704 4156 11756 4208
rect 13728 4156 13780 4208
rect 6368 4131 6420 4140
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 10324 4088 10376 4140
rect 3056 4020 3108 4072
rect 5816 4020 5868 4072
rect 10600 4063 10652 4072
rect 10600 4029 10609 4063
rect 10609 4029 10643 4063
rect 10643 4029 10652 4063
rect 10600 4020 10652 4029
rect 14372 4020 14424 4072
rect 2780 3884 2832 3936
rect 8024 3884 8076 3936
rect 12900 3884 12952 3936
rect 4424 3782 4476 3834
rect 4488 3782 4540 3834
rect 4552 3782 4604 3834
rect 4616 3782 4668 3834
rect 4680 3782 4732 3834
rect 11372 3782 11424 3834
rect 11436 3782 11488 3834
rect 11500 3782 11552 3834
rect 11564 3782 11616 3834
rect 11628 3782 11680 3834
rect 18320 3782 18372 3834
rect 18384 3782 18436 3834
rect 18448 3782 18500 3834
rect 18512 3782 18564 3834
rect 18576 3782 18628 3834
rect 25268 3782 25320 3834
rect 25332 3782 25384 3834
rect 25396 3782 25448 3834
rect 25460 3782 25512 3834
rect 25524 3782 25576 3834
rect 20 3680 72 3732
rect 6092 3680 6144 3732
rect 3056 3655 3108 3664
rect 3056 3621 3065 3655
rect 3065 3621 3099 3655
rect 3099 3621 3108 3655
rect 3056 3612 3108 3621
rect 7472 3612 7524 3664
rect 2780 3544 2832 3596
rect 2044 3476 2096 3528
rect 10324 3544 10376 3596
rect 16120 3723 16172 3732
rect 16120 3689 16129 3723
rect 16129 3689 16163 3723
rect 16163 3689 16172 3723
rect 16120 3680 16172 3689
rect 14004 3612 14056 3664
rect 3976 3408 4028 3460
rect 4252 3451 4304 3460
rect 4252 3417 4261 3451
rect 4261 3417 4295 3451
rect 4295 3417 4304 3451
rect 4252 3408 4304 3417
rect 8484 3476 8536 3528
rect 11980 3476 12032 3528
rect 16212 3519 16264 3528
rect 16212 3485 16221 3519
rect 16221 3485 16255 3519
rect 16255 3485 16264 3519
rect 16212 3476 16264 3485
rect 6368 3408 6420 3460
rect 6552 3408 6604 3460
rect 10600 3408 10652 3460
rect 10784 3408 10836 3460
rect 14464 3408 14516 3460
rect 4896 3340 4948 3392
rect 7748 3340 7800 3392
rect 8024 3340 8076 3392
rect 7898 3238 7950 3290
rect 7962 3238 8014 3290
rect 8026 3238 8078 3290
rect 8090 3238 8142 3290
rect 8154 3238 8206 3290
rect 14846 3238 14898 3290
rect 14910 3238 14962 3290
rect 14974 3238 15026 3290
rect 15038 3238 15090 3290
rect 15102 3238 15154 3290
rect 21794 3238 21846 3290
rect 21858 3238 21910 3290
rect 21922 3238 21974 3290
rect 21986 3238 22038 3290
rect 22050 3238 22102 3290
rect 2780 3111 2832 3120
rect 2780 3077 2789 3111
rect 2789 3077 2823 3111
rect 2823 3077 2832 3111
rect 2780 3068 2832 3077
rect 4344 3111 4396 3120
rect 4344 3077 4353 3111
rect 4353 3077 4387 3111
rect 4387 3077 4396 3111
rect 4344 3068 4396 3077
rect 4252 3000 4304 3052
rect 5816 3043 5868 3052
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 5816 3000 5868 3009
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 10324 3136 10376 3188
rect 10600 3136 10652 3188
rect 14464 3179 14516 3188
rect 8484 3111 8536 3120
rect 8484 3077 8493 3111
rect 8493 3077 8527 3111
rect 8527 3077 8536 3111
rect 8484 3068 8536 3077
rect 10968 3068 11020 3120
rect 14464 3145 14473 3179
rect 14473 3145 14507 3179
rect 14507 3145 14516 3179
rect 14464 3136 14516 3145
rect 10784 3043 10836 3052
rect 10784 3009 10793 3043
rect 10793 3009 10827 3043
rect 10827 3009 10836 3043
rect 10784 3000 10836 3009
rect 7748 2932 7800 2984
rect 11980 2932 12032 2984
rect 14740 3000 14792 3052
rect 4424 2694 4476 2746
rect 4488 2694 4540 2746
rect 4552 2694 4604 2746
rect 4616 2694 4668 2746
rect 4680 2694 4732 2746
rect 11372 2694 11424 2746
rect 11436 2694 11488 2746
rect 11500 2694 11552 2746
rect 11564 2694 11616 2746
rect 11628 2694 11680 2746
rect 18320 2694 18372 2746
rect 18384 2694 18436 2746
rect 18448 2694 18500 2746
rect 18512 2694 18564 2746
rect 18576 2694 18628 2746
rect 25268 2694 25320 2746
rect 25332 2694 25384 2746
rect 25396 2694 25448 2746
rect 25460 2694 25512 2746
rect 25524 2694 25576 2746
rect 5264 2592 5316 2644
rect 23296 2567 23348 2576
rect 23296 2533 23305 2567
rect 23305 2533 23339 2567
rect 23339 2533 23348 2567
rect 23296 2524 23348 2533
rect 2780 2456 2832 2508
rect 2044 2320 2096 2372
rect 16396 2320 16448 2372
rect 23204 2320 23256 2372
rect 7898 2150 7950 2202
rect 7962 2150 8014 2202
rect 8026 2150 8078 2202
rect 8090 2150 8142 2202
rect 8154 2150 8206 2202
rect 14846 2150 14898 2202
rect 14910 2150 14962 2202
rect 14974 2150 15026 2202
rect 15038 2150 15090 2202
rect 15102 2150 15154 2202
rect 21794 2150 21846 2202
rect 21858 2150 21910 2202
rect 21922 2150 21974 2202
rect 21986 2150 22038 2202
rect 22050 2150 22102 2202
<< metal2 >>
rect 18050 29200 18106 30000
rect 4424 27772 4732 27781
rect 4424 27770 4430 27772
rect 4486 27770 4510 27772
rect 4566 27770 4590 27772
rect 4646 27770 4670 27772
rect 4726 27770 4732 27772
rect 4486 27718 4488 27770
rect 4668 27718 4670 27770
rect 4424 27716 4430 27718
rect 4486 27716 4510 27718
rect 4566 27716 4590 27718
rect 4646 27716 4670 27718
rect 4726 27716 4732 27718
rect 4424 27707 4732 27716
rect 11372 27772 11680 27781
rect 11372 27770 11378 27772
rect 11434 27770 11458 27772
rect 11514 27770 11538 27772
rect 11594 27770 11618 27772
rect 11674 27770 11680 27772
rect 11434 27718 11436 27770
rect 11616 27718 11618 27770
rect 11372 27716 11378 27718
rect 11434 27716 11458 27718
rect 11514 27716 11538 27718
rect 11594 27716 11618 27718
rect 11674 27716 11680 27718
rect 11372 27707 11680 27716
rect 18064 27606 18092 29200
rect 18320 27772 18628 27781
rect 18320 27770 18326 27772
rect 18382 27770 18406 27772
rect 18462 27770 18486 27772
rect 18542 27770 18566 27772
rect 18622 27770 18628 27772
rect 18382 27718 18384 27770
rect 18564 27718 18566 27770
rect 18320 27716 18326 27718
rect 18382 27716 18406 27718
rect 18462 27716 18486 27718
rect 18542 27716 18566 27718
rect 18622 27716 18628 27718
rect 18320 27707 18628 27716
rect 25268 27772 25576 27781
rect 25268 27770 25274 27772
rect 25330 27770 25354 27772
rect 25410 27770 25434 27772
rect 25490 27770 25514 27772
rect 25570 27770 25576 27772
rect 25330 27718 25332 27770
rect 25512 27718 25514 27770
rect 25268 27716 25274 27718
rect 25330 27716 25354 27718
rect 25410 27716 25434 27718
rect 25490 27716 25514 27718
rect 25570 27716 25576 27718
rect 25268 27707 25576 27716
rect 18052 27600 18104 27606
rect 18052 27542 18104 27548
rect 18144 27328 18196 27334
rect 18144 27270 18196 27276
rect 7898 27228 8206 27237
rect 7898 27226 7904 27228
rect 7960 27226 7984 27228
rect 8040 27226 8064 27228
rect 8120 27226 8144 27228
rect 8200 27226 8206 27228
rect 7960 27174 7962 27226
rect 8142 27174 8144 27226
rect 7898 27172 7904 27174
rect 7960 27172 7984 27174
rect 8040 27172 8064 27174
rect 8120 27172 8144 27174
rect 8200 27172 8206 27174
rect 7898 27163 8206 27172
rect 14846 27228 15154 27237
rect 14846 27226 14852 27228
rect 14908 27226 14932 27228
rect 14988 27226 15012 27228
rect 15068 27226 15092 27228
rect 15148 27226 15154 27228
rect 14908 27174 14910 27226
rect 15090 27174 15092 27226
rect 14846 27172 14852 27174
rect 14908 27172 14932 27174
rect 14988 27172 15012 27174
rect 15068 27172 15092 27174
rect 15148 27172 15154 27174
rect 14846 27163 15154 27172
rect 4424 26684 4732 26693
rect 4424 26682 4430 26684
rect 4486 26682 4510 26684
rect 4566 26682 4590 26684
rect 4646 26682 4670 26684
rect 4726 26682 4732 26684
rect 4486 26630 4488 26682
rect 4668 26630 4670 26682
rect 4424 26628 4430 26630
rect 4486 26628 4510 26630
rect 4566 26628 4590 26630
rect 4646 26628 4670 26630
rect 4726 26628 4732 26630
rect 4424 26619 4732 26628
rect 11372 26684 11680 26693
rect 11372 26682 11378 26684
rect 11434 26682 11458 26684
rect 11514 26682 11538 26684
rect 11594 26682 11618 26684
rect 11674 26682 11680 26684
rect 11434 26630 11436 26682
rect 11616 26630 11618 26682
rect 11372 26628 11378 26630
rect 11434 26628 11458 26630
rect 11514 26628 11538 26630
rect 11594 26628 11618 26630
rect 11674 26628 11680 26630
rect 11372 26619 11680 26628
rect 7898 26140 8206 26149
rect 7898 26138 7904 26140
rect 7960 26138 7984 26140
rect 8040 26138 8064 26140
rect 8120 26138 8144 26140
rect 8200 26138 8206 26140
rect 7960 26086 7962 26138
rect 8142 26086 8144 26138
rect 7898 26084 7904 26086
rect 7960 26084 7984 26086
rect 8040 26084 8064 26086
rect 8120 26084 8144 26086
rect 8200 26084 8206 26086
rect 7898 26075 8206 26084
rect 14846 26140 15154 26149
rect 14846 26138 14852 26140
rect 14908 26138 14932 26140
rect 14988 26138 15012 26140
rect 15068 26138 15092 26140
rect 15148 26138 15154 26140
rect 14908 26086 14910 26138
rect 15090 26086 15092 26138
rect 14846 26084 14852 26086
rect 14908 26084 14932 26086
rect 14988 26084 15012 26086
rect 15068 26084 15092 26086
rect 15148 26084 15154 26086
rect 14846 26075 15154 26084
rect 4424 25596 4732 25605
rect 4424 25594 4430 25596
rect 4486 25594 4510 25596
rect 4566 25594 4590 25596
rect 4646 25594 4670 25596
rect 4726 25594 4732 25596
rect 4486 25542 4488 25594
rect 4668 25542 4670 25594
rect 4424 25540 4430 25542
rect 4486 25540 4510 25542
rect 4566 25540 4590 25542
rect 4646 25540 4670 25542
rect 4726 25540 4732 25542
rect 4424 25531 4732 25540
rect 11372 25596 11680 25605
rect 11372 25594 11378 25596
rect 11434 25594 11458 25596
rect 11514 25594 11538 25596
rect 11594 25594 11618 25596
rect 11674 25594 11680 25596
rect 11434 25542 11436 25594
rect 11616 25542 11618 25594
rect 11372 25540 11378 25542
rect 11434 25540 11458 25542
rect 11514 25540 11538 25542
rect 11594 25540 11618 25542
rect 11674 25540 11680 25542
rect 11372 25531 11680 25540
rect 7898 25052 8206 25061
rect 7898 25050 7904 25052
rect 7960 25050 7984 25052
rect 8040 25050 8064 25052
rect 8120 25050 8144 25052
rect 8200 25050 8206 25052
rect 7960 24998 7962 25050
rect 8142 24998 8144 25050
rect 7898 24996 7904 24998
rect 7960 24996 7984 24998
rect 8040 24996 8064 24998
rect 8120 24996 8144 24998
rect 8200 24996 8206 24998
rect 7898 24987 8206 24996
rect 14846 25052 15154 25061
rect 14846 25050 14852 25052
rect 14908 25050 14932 25052
rect 14988 25050 15012 25052
rect 15068 25050 15092 25052
rect 15148 25050 15154 25052
rect 14908 24998 14910 25050
rect 15090 24998 15092 25050
rect 14846 24996 14852 24998
rect 14908 24996 14932 24998
rect 14988 24996 15012 24998
rect 15068 24996 15092 24998
rect 15148 24996 15154 24998
rect 14846 24987 15154 24996
rect 6368 24812 6420 24818
rect 6368 24754 6420 24760
rect 1492 24608 1544 24614
rect 1490 24576 1492 24585
rect 1544 24576 1546 24585
rect 1490 24511 1546 24520
rect 4424 24508 4732 24517
rect 4424 24506 4430 24508
rect 4486 24506 4510 24508
rect 4566 24506 4590 24508
rect 4646 24506 4670 24508
rect 4726 24506 4732 24508
rect 4486 24454 4488 24506
rect 4668 24454 4670 24506
rect 4424 24452 4430 24454
rect 4486 24452 4510 24454
rect 4566 24452 4590 24454
rect 4646 24452 4670 24454
rect 4726 24452 4732 24454
rect 4424 24443 4732 24452
rect 4424 23420 4732 23429
rect 4424 23418 4430 23420
rect 4486 23418 4510 23420
rect 4566 23418 4590 23420
rect 4646 23418 4670 23420
rect 4726 23418 4732 23420
rect 4486 23366 4488 23418
rect 4668 23366 4670 23418
rect 4424 23364 4430 23366
rect 4486 23364 4510 23366
rect 4566 23364 4590 23366
rect 4646 23364 4670 23366
rect 4726 23364 4732 23366
rect 4424 23355 4732 23364
rect 4424 22332 4732 22341
rect 4424 22330 4430 22332
rect 4486 22330 4510 22332
rect 4566 22330 4590 22332
rect 4646 22330 4670 22332
rect 4726 22330 4732 22332
rect 4486 22278 4488 22330
rect 4668 22278 4670 22330
rect 4424 22276 4430 22278
rect 4486 22276 4510 22278
rect 4566 22276 4590 22278
rect 4646 22276 4670 22278
rect 4726 22276 4732 22278
rect 4424 22267 4732 22276
rect 4424 21244 4732 21253
rect 4424 21242 4430 21244
rect 4486 21242 4510 21244
rect 4566 21242 4590 21244
rect 4646 21242 4670 21244
rect 4726 21242 4732 21244
rect 4486 21190 4488 21242
rect 4668 21190 4670 21242
rect 4424 21188 4430 21190
rect 4486 21188 4510 21190
rect 4566 21188 4590 21190
rect 4646 21188 4670 21190
rect 4726 21188 4732 21190
rect 4424 21179 4732 21188
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3988 20262 4016 20402
rect 3792 20256 3844 20262
rect 3792 20198 3844 20204
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3160 16574 3188 19790
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3068 16546 3188 16574
rect 2964 16516 3016 16522
rect 2964 16458 3016 16464
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1688 13326 1716 13806
rect 1964 13802 1992 14962
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 1952 13796 2004 13802
rect 1952 13738 2004 13744
rect 1964 13530 1992 13738
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1504 10810 1532 11086
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1780 10130 1808 13126
rect 1768 10124 1820 10130
rect 1768 10066 1820 10072
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1504 9518 1532 9998
rect 2056 9654 2084 14758
rect 2136 14272 2188 14278
rect 2136 14214 2188 14220
rect 2148 10742 2176 14214
rect 2424 12714 2452 14962
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2688 14340 2740 14346
rect 2688 14282 2740 14288
rect 2700 13394 2728 14282
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2700 12986 2728 13330
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2412 12708 2464 12714
rect 2412 12650 2464 12656
rect 2792 11218 2820 14214
rect 2884 13938 2912 14486
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2884 13258 2912 13874
rect 2976 13802 3004 16458
rect 2964 13796 3016 13802
rect 2964 13738 3016 13744
rect 2872 13252 2924 13258
rect 2872 13194 2924 13200
rect 2884 12918 2912 13194
rect 2976 13190 3004 13738
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2976 12850 3004 13126
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2136 10736 2188 10742
rect 2136 10678 2188 10684
rect 2044 9648 2096 9654
rect 2044 9590 2096 9596
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1768 7812 1820 7818
rect 1768 7754 1820 7760
rect 1780 7410 1808 7754
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 3068 6914 3096 16546
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3252 14074 3280 14350
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 3148 14000 3200 14006
rect 3148 13942 3200 13948
rect 3160 13394 3188 13942
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 3160 11354 3188 13330
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 3252 10266 3280 13806
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 3344 9518 3372 12786
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 9042 3280 9318
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 3252 8498 3280 8978
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3252 7954 3280 8434
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3252 7546 3280 7890
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3068 6886 3188 6914
rect 3160 6798 3188 6886
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 2332 6390 2360 6734
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2320 6384 2372 6390
rect 2320 6326 2372 6332
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2792 5166 2820 6054
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1780 4554 1808 4966
rect 2792 4690 2820 5102
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 1768 4548 1820 4554
rect 1768 4490 1820 4496
rect 2792 3942 2820 4626
rect 3068 4554 3096 6598
rect 3436 6322 3464 19654
rect 3804 16574 3832 20198
rect 3988 19854 4016 20198
rect 4424 20156 4732 20165
rect 4424 20154 4430 20156
rect 4486 20154 4510 20156
rect 4566 20154 4590 20156
rect 4646 20154 4670 20156
rect 4726 20154 4732 20156
rect 4486 20102 4488 20154
rect 4668 20102 4670 20154
rect 4424 20100 4430 20102
rect 4486 20100 4510 20102
rect 4566 20100 4590 20102
rect 4646 20100 4670 20102
rect 4726 20100 4732 20102
rect 4424 20091 4732 20100
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 4424 19068 4732 19077
rect 4424 19066 4430 19068
rect 4486 19066 4510 19068
rect 4566 19066 4590 19068
rect 4646 19066 4670 19068
rect 4726 19066 4732 19068
rect 4486 19014 4488 19066
rect 4668 19014 4670 19066
rect 4424 19012 4430 19014
rect 4486 19012 4510 19014
rect 4566 19012 4590 19014
rect 4646 19012 4670 19014
rect 4726 19012 4732 19014
rect 4424 19003 4732 19012
rect 4424 17980 4732 17989
rect 4424 17978 4430 17980
rect 4486 17978 4510 17980
rect 4566 17978 4590 17980
rect 4646 17978 4670 17980
rect 4726 17978 4732 17980
rect 4486 17926 4488 17978
rect 4668 17926 4670 17978
rect 4424 17924 4430 17926
rect 4486 17924 4510 17926
rect 4566 17924 4590 17926
rect 4646 17924 4670 17926
rect 4726 17924 4732 17926
rect 4424 17915 4732 17924
rect 5632 17264 5684 17270
rect 5632 17206 5684 17212
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4424 16892 4732 16901
rect 4424 16890 4430 16892
rect 4486 16890 4510 16892
rect 4566 16890 4590 16892
rect 4646 16890 4670 16892
rect 4726 16890 4732 16892
rect 4486 16838 4488 16890
rect 4668 16838 4670 16890
rect 4424 16836 4430 16838
rect 4486 16836 4510 16838
rect 4566 16836 4590 16838
rect 4646 16836 4670 16838
rect 4726 16836 4732 16838
rect 4424 16827 4732 16836
rect 4816 16590 4844 16934
rect 3712 16546 3832 16574
rect 4804 16584 4856 16590
rect 3608 14952 3660 14958
rect 3608 14894 3660 14900
rect 3620 13870 3648 14894
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3528 9994 3556 12718
rect 3516 9988 3568 9994
rect 3516 9930 3568 9936
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3528 8090 3556 8366
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3712 7818 3740 16546
rect 4804 16526 4856 16532
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3804 14550 3832 15982
rect 3792 14544 3844 14550
rect 3792 14486 3844 14492
rect 3804 14414 3832 14486
rect 4080 14414 4108 16390
rect 4908 16250 4936 17138
rect 4988 17060 5040 17066
rect 4988 17002 5040 17008
rect 5000 16590 5028 17002
rect 5644 16658 5672 17206
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 4896 16244 4948 16250
rect 4896 16186 4948 16192
rect 5552 16182 5580 16390
rect 5540 16176 5592 16182
rect 5540 16118 5592 16124
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 4172 15026 4200 15982
rect 4424 15804 4732 15813
rect 4424 15802 4430 15804
rect 4486 15802 4510 15804
rect 4566 15802 4590 15804
rect 4646 15802 4670 15804
rect 4726 15802 4732 15804
rect 4486 15750 4488 15802
rect 4668 15750 4670 15802
rect 4424 15748 4430 15750
rect 4486 15748 4510 15750
rect 4566 15748 4590 15750
rect 4646 15748 4670 15750
rect 4726 15748 4732 15750
rect 4424 15739 4732 15748
rect 4908 15162 4936 16050
rect 5000 15570 5028 16050
rect 4988 15564 5040 15570
rect 4988 15506 5040 15512
rect 5460 15366 5488 16050
rect 5644 15706 5672 16594
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 5736 16454 5764 16526
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5736 16114 5764 16390
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5644 15366 5672 15642
rect 5736 15502 5764 16050
rect 6380 15978 6408 24754
rect 11372 24508 11680 24517
rect 11372 24506 11378 24508
rect 11434 24506 11458 24508
rect 11514 24506 11538 24508
rect 11594 24506 11618 24508
rect 11674 24506 11680 24508
rect 11434 24454 11436 24506
rect 11616 24454 11618 24506
rect 11372 24452 11378 24454
rect 11434 24452 11458 24454
rect 11514 24452 11538 24454
rect 11594 24452 11618 24454
rect 11674 24452 11680 24454
rect 11372 24443 11680 24452
rect 7898 23964 8206 23973
rect 7898 23962 7904 23964
rect 7960 23962 7984 23964
rect 8040 23962 8064 23964
rect 8120 23962 8144 23964
rect 8200 23962 8206 23964
rect 7960 23910 7962 23962
rect 8142 23910 8144 23962
rect 7898 23908 7904 23910
rect 7960 23908 7984 23910
rect 8040 23908 8064 23910
rect 8120 23908 8144 23910
rect 8200 23908 8206 23910
rect 7898 23899 8206 23908
rect 14846 23964 15154 23973
rect 14846 23962 14852 23964
rect 14908 23962 14932 23964
rect 14988 23962 15012 23964
rect 15068 23962 15092 23964
rect 15148 23962 15154 23964
rect 14908 23910 14910 23962
rect 15090 23910 15092 23962
rect 14846 23908 14852 23910
rect 14908 23908 14932 23910
rect 14988 23908 15012 23910
rect 15068 23908 15092 23910
rect 15148 23908 15154 23910
rect 14846 23899 15154 23908
rect 11372 23420 11680 23429
rect 11372 23418 11378 23420
rect 11434 23418 11458 23420
rect 11514 23418 11538 23420
rect 11594 23418 11618 23420
rect 11674 23418 11680 23420
rect 11434 23366 11436 23418
rect 11616 23366 11618 23418
rect 11372 23364 11378 23366
rect 11434 23364 11458 23366
rect 11514 23364 11538 23366
rect 11594 23364 11618 23366
rect 11674 23364 11680 23366
rect 11372 23355 11680 23364
rect 7898 22876 8206 22885
rect 7898 22874 7904 22876
rect 7960 22874 7984 22876
rect 8040 22874 8064 22876
rect 8120 22874 8144 22876
rect 8200 22874 8206 22876
rect 7960 22822 7962 22874
rect 8142 22822 8144 22874
rect 7898 22820 7904 22822
rect 7960 22820 7984 22822
rect 8040 22820 8064 22822
rect 8120 22820 8144 22822
rect 8200 22820 8206 22822
rect 7898 22811 8206 22820
rect 14846 22876 15154 22885
rect 14846 22874 14852 22876
rect 14908 22874 14932 22876
rect 14988 22874 15012 22876
rect 15068 22874 15092 22876
rect 15148 22874 15154 22876
rect 14908 22822 14910 22874
rect 15090 22822 15092 22874
rect 14846 22820 14852 22822
rect 14908 22820 14932 22822
rect 14988 22820 15012 22822
rect 15068 22820 15092 22822
rect 15148 22820 15154 22822
rect 14846 22811 15154 22820
rect 11372 22332 11680 22341
rect 11372 22330 11378 22332
rect 11434 22330 11458 22332
rect 11514 22330 11538 22332
rect 11594 22330 11618 22332
rect 11674 22330 11680 22332
rect 11434 22278 11436 22330
rect 11616 22278 11618 22330
rect 11372 22276 11378 22278
rect 11434 22276 11458 22278
rect 11514 22276 11538 22278
rect 11594 22276 11618 22278
rect 11674 22276 11680 22278
rect 11372 22267 11680 22276
rect 7898 21788 8206 21797
rect 7898 21786 7904 21788
rect 7960 21786 7984 21788
rect 8040 21786 8064 21788
rect 8120 21786 8144 21788
rect 8200 21786 8206 21788
rect 7960 21734 7962 21786
rect 8142 21734 8144 21786
rect 7898 21732 7904 21734
rect 7960 21732 7984 21734
rect 8040 21732 8064 21734
rect 8120 21732 8144 21734
rect 8200 21732 8206 21734
rect 7898 21723 8206 21732
rect 14846 21788 15154 21797
rect 14846 21786 14852 21788
rect 14908 21786 14932 21788
rect 14988 21786 15012 21788
rect 15068 21786 15092 21788
rect 15148 21786 15154 21788
rect 14908 21734 14910 21786
rect 15090 21734 15092 21786
rect 14846 21732 14852 21734
rect 14908 21732 14932 21734
rect 14988 21732 15012 21734
rect 15068 21732 15092 21734
rect 15148 21732 15154 21734
rect 14846 21723 15154 21732
rect 11372 21244 11680 21253
rect 11372 21242 11378 21244
rect 11434 21242 11458 21244
rect 11514 21242 11538 21244
rect 11594 21242 11618 21244
rect 11674 21242 11680 21244
rect 11434 21190 11436 21242
rect 11616 21190 11618 21242
rect 11372 21188 11378 21190
rect 11434 21188 11458 21190
rect 11514 21188 11538 21190
rect 11594 21188 11618 21190
rect 11674 21188 11680 21190
rect 11372 21179 11680 21188
rect 7898 20700 8206 20709
rect 7898 20698 7904 20700
rect 7960 20698 7984 20700
rect 8040 20698 8064 20700
rect 8120 20698 8144 20700
rect 8200 20698 8206 20700
rect 7960 20646 7962 20698
rect 8142 20646 8144 20698
rect 7898 20644 7904 20646
rect 7960 20644 7984 20646
rect 8040 20644 8064 20646
rect 8120 20644 8144 20646
rect 8200 20644 8206 20646
rect 7898 20635 8206 20644
rect 14846 20700 15154 20709
rect 14846 20698 14852 20700
rect 14908 20698 14932 20700
rect 14988 20698 15012 20700
rect 15068 20698 15092 20700
rect 15148 20698 15154 20700
rect 14908 20646 14910 20698
rect 15090 20646 15092 20698
rect 14846 20644 14852 20646
rect 14908 20644 14932 20646
rect 14988 20644 15012 20646
rect 15068 20644 15092 20646
rect 15148 20644 15154 20646
rect 14846 20635 15154 20644
rect 11372 20156 11680 20165
rect 11372 20154 11378 20156
rect 11434 20154 11458 20156
rect 11514 20154 11538 20156
rect 11594 20154 11618 20156
rect 11674 20154 11680 20156
rect 11434 20102 11436 20154
rect 11616 20102 11618 20154
rect 11372 20100 11378 20102
rect 11434 20100 11458 20102
rect 11514 20100 11538 20102
rect 11594 20100 11618 20102
rect 11674 20100 11680 20102
rect 11372 20091 11680 20100
rect 7898 19612 8206 19621
rect 7898 19610 7904 19612
rect 7960 19610 7984 19612
rect 8040 19610 8064 19612
rect 8120 19610 8144 19612
rect 8200 19610 8206 19612
rect 7960 19558 7962 19610
rect 8142 19558 8144 19610
rect 7898 19556 7904 19558
rect 7960 19556 7984 19558
rect 8040 19556 8064 19558
rect 8120 19556 8144 19558
rect 8200 19556 8206 19558
rect 7898 19547 8206 19556
rect 14846 19612 15154 19621
rect 14846 19610 14852 19612
rect 14908 19610 14932 19612
rect 14988 19610 15012 19612
rect 15068 19610 15092 19612
rect 15148 19610 15154 19612
rect 14908 19558 14910 19610
rect 15090 19558 15092 19610
rect 14846 19556 14852 19558
rect 14908 19556 14932 19558
rect 14988 19556 15012 19558
rect 15068 19556 15092 19558
rect 15148 19556 15154 19558
rect 14846 19547 15154 19556
rect 11372 19068 11680 19077
rect 11372 19066 11378 19068
rect 11434 19066 11458 19068
rect 11514 19066 11538 19068
rect 11594 19066 11618 19068
rect 11674 19066 11680 19068
rect 11434 19014 11436 19066
rect 11616 19014 11618 19066
rect 11372 19012 11378 19014
rect 11434 19012 11458 19014
rect 11514 19012 11538 19014
rect 11594 19012 11618 19014
rect 11674 19012 11680 19014
rect 11372 19003 11680 19012
rect 7898 18524 8206 18533
rect 7898 18522 7904 18524
rect 7960 18522 7984 18524
rect 8040 18522 8064 18524
rect 8120 18522 8144 18524
rect 8200 18522 8206 18524
rect 7960 18470 7962 18522
rect 8142 18470 8144 18522
rect 7898 18468 7904 18470
rect 7960 18468 7984 18470
rect 8040 18468 8064 18470
rect 8120 18468 8144 18470
rect 8200 18468 8206 18470
rect 7898 18459 8206 18468
rect 14846 18524 15154 18533
rect 14846 18522 14852 18524
rect 14908 18522 14932 18524
rect 14988 18522 15012 18524
rect 15068 18522 15092 18524
rect 15148 18522 15154 18524
rect 14908 18470 14910 18522
rect 15090 18470 15092 18522
rect 14846 18468 14852 18470
rect 14908 18468 14932 18470
rect 14988 18468 15012 18470
rect 15068 18468 15092 18470
rect 15148 18468 15154 18470
rect 14846 18459 15154 18468
rect 11372 17980 11680 17989
rect 11372 17978 11378 17980
rect 11434 17978 11458 17980
rect 11514 17978 11538 17980
rect 11594 17978 11618 17980
rect 11674 17978 11680 17980
rect 11434 17926 11436 17978
rect 11616 17926 11618 17978
rect 11372 17924 11378 17926
rect 11434 17924 11458 17926
rect 11514 17924 11538 17926
rect 11594 17924 11618 17926
rect 11674 17924 11680 17926
rect 11372 17915 11680 17924
rect 7898 17436 8206 17445
rect 7898 17434 7904 17436
rect 7960 17434 7984 17436
rect 8040 17434 8064 17436
rect 8120 17434 8144 17436
rect 8200 17434 8206 17436
rect 7960 17382 7962 17434
rect 8142 17382 8144 17434
rect 7898 17380 7904 17382
rect 7960 17380 7984 17382
rect 8040 17380 8064 17382
rect 8120 17380 8144 17382
rect 8200 17380 8206 17382
rect 7898 17371 8206 17380
rect 14846 17436 15154 17445
rect 14846 17434 14852 17436
rect 14908 17434 14932 17436
rect 14988 17434 15012 17436
rect 15068 17434 15092 17436
rect 15148 17434 15154 17436
rect 14908 17382 14910 17434
rect 15090 17382 15092 17434
rect 14846 17380 14852 17382
rect 14908 17380 14932 17382
rect 14988 17380 15012 17382
rect 15068 17380 15092 17382
rect 15148 17380 15154 17382
rect 14846 17371 15154 17380
rect 7564 17264 7616 17270
rect 7564 17206 7616 17212
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7392 16574 7420 17002
rect 7576 16658 7604 17206
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7024 16546 7420 16574
rect 6644 16516 6696 16522
rect 6644 16458 6696 16464
rect 6656 16114 6684 16458
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6368 15972 6420 15978
rect 6368 15914 6420 15920
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 6368 15496 6420 15502
rect 6368 15438 6420 15444
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5460 15162 5488 15302
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3976 14272 4028 14278
rect 3976 14214 4028 14220
rect 3896 13938 3924 14214
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3896 10742 3924 12650
rect 3988 11286 4016 14214
rect 4080 14006 4108 14350
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3988 10810 4016 11086
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3884 10736 3936 10742
rect 3884 10678 3936 10684
rect 3988 10690 4016 10746
rect 3988 10662 4108 10690
rect 4080 10606 4108 10662
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4080 9042 4108 10542
rect 4172 10470 4200 14962
rect 4424 14716 4732 14725
rect 4424 14714 4430 14716
rect 4486 14714 4510 14716
rect 4566 14714 4590 14716
rect 4646 14714 4670 14716
rect 4726 14714 4732 14716
rect 4486 14662 4488 14714
rect 4668 14662 4670 14714
rect 4424 14660 4430 14662
rect 4486 14660 4510 14662
rect 4566 14660 4590 14662
rect 4646 14660 4670 14662
rect 4726 14660 4732 14662
rect 4424 14651 4732 14660
rect 5080 14408 5132 14414
rect 5080 14350 5132 14356
rect 4424 13628 4732 13637
rect 4424 13626 4430 13628
rect 4486 13626 4510 13628
rect 4566 13626 4590 13628
rect 4646 13626 4670 13628
rect 4726 13626 4732 13628
rect 4486 13574 4488 13626
rect 4668 13574 4670 13626
rect 4424 13572 4430 13574
rect 4486 13572 4510 13574
rect 4566 13572 4590 13574
rect 4646 13572 4670 13574
rect 4726 13572 4732 13574
rect 4424 13563 4732 13572
rect 5092 13326 5120 14350
rect 5816 13796 5868 13802
rect 5816 13738 5868 13744
rect 5080 13320 5132 13326
rect 4250 13288 4306 13297
rect 5080 13262 5132 13268
rect 4250 13223 4252 13232
rect 4304 13223 4306 13232
rect 4252 13194 4304 13200
rect 4264 12986 4292 13194
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4424 12540 4732 12549
rect 4424 12538 4430 12540
rect 4486 12538 4510 12540
rect 4566 12538 4590 12540
rect 4646 12538 4670 12540
rect 4726 12538 4732 12540
rect 4486 12486 4488 12538
rect 4668 12486 4670 12538
rect 4424 12484 4430 12486
rect 4486 12484 4510 12486
rect 4566 12484 4590 12486
rect 4646 12484 4670 12486
rect 4726 12484 4732 12486
rect 4424 12475 4732 12484
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4264 11218 4292 12038
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4356 10742 4384 11494
rect 4424 11452 4732 11461
rect 4424 11450 4430 11452
rect 4486 11450 4510 11452
rect 4566 11450 4590 11452
rect 4646 11450 4670 11452
rect 4726 11450 4732 11452
rect 4486 11398 4488 11450
rect 4668 11398 4670 11450
rect 4424 11396 4430 11398
rect 4486 11396 4510 11398
rect 4566 11396 4590 11398
rect 4646 11396 4670 11398
rect 4726 11396 4732 11398
rect 4424 11387 4732 11396
rect 4816 11082 4844 12582
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4424 10364 4732 10373
rect 4424 10362 4430 10364
rect 4486 10362 4510 10364
rect 4566 10362 4590 10364
rect 4646 10362 4670 10364
rect 4726 10362 4732 10364
rect 4486 10310 4488 10362
rect 4668 10310 4670 10362
rect 4424 10308 4430 10310
rect 4486 10308 4510 10310
rect 4566 10308 4590 10310
rect 4646 10308 4670 10310
rect 4726 10308 4732 10310
rect 4424 10299 4732 10308
rect 5000 9654 5028 13126
rect 5092 12850 5120 13262
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5460 10674 5488 13126
rect 5828 10674 5856 13738
rect 6380 13394 6408 15438
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 6564 14482 6592 14962
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6460 14272 6512 14278
rect 6460 14214 6512 14220
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6196 12238 6224 13126
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6380 11354 6408 13330
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5828 10266 5856 10406
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 6380 10130 6408 10542
rect 6472 10130 6500 14214
rect 6656 14006 6684 15438
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6564 13190 6592 13874
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 4424 9276 4732 9285
rect 4424 9274 4430 9276
rect 4486 9274 4510 9276
rect 4566 9274 4590 9276
rect 4646 9274 4670 9276
rect 4726 9274 4732 9276
rect 4486 9222 4488 9274
rect 4668 9222 4670 9274
rect 4424 9220 4430 9222
rect 4486 9220 4510 9222
rect 4566 9220 4590 9222
rect 4646 9220 4670 9222
rect 4726 9220 4732 9222
rect 4424 9211 4732 9220
rect 6380 9042 6408 10066
rect 6564 9518 6592 13126
rect 6656 10606 6684 13942
rect 6748 13870 6776 15506
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6828 13796 6880 13802
rect 6828 13738 6880 13744
rect 6840 13394 6868 13738
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6932 9994 6960 12582
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 7024 9042 7052 16546
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7208 14414 7236 15846
rect 7392 15706 7420 16050
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7380 15496 7432 15502
rect 7484 15484 7512 15982
rect 7432 15456 7512 15484
rect 7380 15438 7432 15444
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7288 14408 7340 14414
rect 7392 14362 7420 15438
rect 7576 14414 7604 16594
rect 7668 16046 7696 16934
rect 7944 16794 7972 17070
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 7760 16250 7788 16594
rect 7898 16348 8206 16357
rect 7898 16346 7904 16348
rect 7960 16346 7984 16348
rect 8040 16346 8064 16348
rect 8120 16346 8144 16348
rect 8200 16346 8206 16348
rect 7960 16294 7962 16346
rect 8142 16294 8144 16346
rect 7898 16292 7904 16294
rect 7960 16292 7984 16294
rect 8040 16292 8064 16294
rect 8120 16292 8144 16294
rect 8200 16292 8206 16294
rect 7898 16283 8206 16292
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 9048 16046 9076 17070
rect 10336 16590 10364 17070
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10428 16726 10456 16934
rect 11372 16892 11680 16901
rect 11372 16890 11378 16892
rect 11434 16890 11458 16892
rect 11514 16890 11538 16892
rect 11594 16890 11618 16892
rect 11674 16890 11680 16892
rect 11434 16838 11436 16890
rect 11616 16838 11618 16890
rect 11372 16836 11378 16838
rect 11434 16836 11458 16838
rect 11514 16836 11538 16838
rect 11594 16836 11618 16838
rect 11674 16836 11680 16838
rect 11372 16827 11680 16836
rect 10416 16720 10468 16726
rect 10416 16662 10468 16668
rect 9312 16584 9364 16590
rect 9588 16584 9640 16590
rect 9312 16526 9364 16532
rect 9508 16532 9588 16538
rect 9508 16526 9640 16532
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 11704 16584 11756 16590
rect 12440 16584 12492 16590
rect 11756 16532 11836 16538
rect 11704 16526 11836 16532
rect 12440 16526 12492 16532
rect 9324 16250 9352 16526
rect 9508 16510 9628 16526
rect 11716 16510 11836 16526
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 8312 15366 8340 15982
rect 9416 15502 9444 15982
rect 9508 15570 9536 16510
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 9496 15564 9548 15570
rect 9496 15506 9548 15512
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 7898 15260 8206 15269
rect 7898 15258 7904 15260
rect 7960 15258 7984 15260
rect 8040 15258 8064 15260
rect 8120 15258 8144 15260
rect 8200 15258 8206 15260
rect 7960 15206 7962 15258
rect 8142 15206 8144 15258
rect 7898 15204 7904 15206
rect 7960 15204 7984 15206
rect 8040 15204 8064 15206
rect 8120 15204 8144 15206
rect 8200 15204 8206 15206
rect 7898 15195 8206 15204
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7340 14356 7420 14362
rect 7288 14350 7420 14356
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7300 14334 7420 14350
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 10742 7328 14214
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 7392 10198 7420 14334
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7484 12850 7512 13670
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7380 10192 7432 10198
rect 7380 10134 7432 10140
rect 7576 9178 7604 14350
rect 7760 14074 7788 14758
rect 7898 14172 8206 14181
rect 7898 14170 7904 14172
rect 7960 14170 7984 14172
rect 8040 14170 8064 14172
rect 8120 14170 8144 14172
rect 8200 14170 8206 14172
rect 7960 14118 7962 14170
rect 8142 14118 8144 14170
rect 7898 14116 7904 14118
rect 7960 14116 7984 14118
rect 8040 14116 8064 14118
rect 8120 14116 8144 14118
rect 8200 14116 8206 14118
rect 7898 14107 8206 14116
rect 8772 14074 8800 15302
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 6656 8922 6684 8978
rect 6564 8906 6684 8922
rect 6552 8900 6684 8906
rect 6604 8894 6684 8900
rect 6552 8842 6604 8848
rect 4804 8560 4856 8566
rect 4804 8502 4856 8508
rect 4424 8188 4732 8197
rect 4424 8186 4430 8188
rect 4486 8186 4510 8188
rect 4566 8186 4590 8188
rect 4646 8186 4670 8188
rect 4726 8186 4732 8188
rect 4486 8134 4488 8186
rect 4668 8134 4670 8186
rect 4424 8132 4430 8134
rect 4486 8132 4510 8134
rect 4566 8132 4590 8134
rect 4646 8132 4670 8134
rect 4726 8132 4732 8134
rect 4424 8123 4732 8132
rect 3700 7812 3752 7818
rect 3700 7754 3752 7760
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4356 7410 4384 7754
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3620 6390 3648 6734
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3804 5914 3832 6054
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3804 4826 3832 5102
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 20 3732 72 3738
rect 20 3674 72 3680
rect 32 800 60 3674
rect 2792 3602 2820 3878
rect 3068 3670 3096 4014
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 2056 2378 2084 3470
rect 2792 3126 2820 3538
rect 4172 3482 4200 4558
rect 3988 3466 4200 3482
rect 3976 3460 4200 3466
rect 4028 3454 4200 3460
rect 4252 3460 4304 3466
rect 3976 3402 4028 3408
rect 4252 3402 4304 3408
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2792 2514 2820 3062
rect 4264 3058 4292 3402
rect 4356 3126 4384 7346
rect 4424 7100 4732 7109
rect 4424 7098 4430 7100
rect 4486 7098 4510 7100
rect 4566 7098 4590 7100
rect 4646 7098 4670 7100
rect 4726 7098 4732 7100
rect 4486 7046 4488 7098
rect 4668 7046 4670 7098
rect 4424 7044 4430 7046
rect 4486 7044 4510 7046
rect 4566 7044 4590 7046
rect 4646 7044 4670 7046
rect 4726 7044 4732 7046
rect 4424 7035 4732 7044
rect 4816 6458 4844 8502
rect 6276 8356 6328 8362
rect 6276 8298 6328 8304
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4424 6012 4732 6021
rect 4424 6010 4430 6012
rect 4486 6010 4510 6012
rect 4566 6010 4590 6012
rect 4646 6010 4670 6012
rect 4726 6010 4732 6012
rect 4486 5958 4488 6010
rect 4668 5958 4670 6010
rect 4424 5956 4430 5958
rect 4486 5956 4510 5958
rect 4566 5956 4590 5958
rect 4646 5956 4670 5958
rect 4726 5956 4732 5958
rect 4424 5947 4732 5956
rect 4908 5030 4936 7686
rect 6196 7478 6224 7686
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5000 7002 5028 7142
rect 5828 7002 5856 7142
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 6196 6914 6224 7414
rect 5906 6896 5962 6905
rect 5906 6831 5962 6840
rect 6104 6886 6224 6914
rect 5920 6662 5948 6831
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5356 6384 5408 6390
rect 5354 6352 5356 6361
rect 5408 6352 5410 6361
rect 5354 6287 5410 6296
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4424 4924 4732 4933
rect 4424 4922 4430 4924
rect 4486 4922 4510 4924
rect 4566 4922 4590 4924
rect 4646 4922 4670 4924
rect 4726 4922 4732 4924
rect 4486 4870 4488 4922
rect 4668 4870 4670 4922
rect 4424 4868 4430 4870
rect 4486 4868 4510 4870
rect 4566 4868 4590 4870
rect 4646 4868 4670 4870
rect 4726 4868 4732 4870
rect 4424 4859 4732 4868
rect 5092 4758 5120 5102
rect 5080 4752 5132 4758
rect 5080 4694 5132 4700
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4632 4214 4660 4422
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 4424 3836 4732 3845
rect 4424 3834 4430 3836
rect 4486 3834 4510 3836
rect 4566 3834 4590 3836
rect 4646 3834 4670 3836
rect 4726 3834 4732 3836
rect 4486 3782 4488 3834
rect 4668 3782 4670 3834
rect 4424 3780 4430 3782
rect 4486 3780 4510 3782
rect 4566 3780 4590 3782
rect 4646 3780 4670 3782
rect 4726 3780 4732 3782
rect 4424 3771 4732 3780
rect 4908 3398 4936 4558
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4424 2748 4732 2757
rect 4424 2746 4430 2748
rect 4486 2746 4510 2748
rect 4566 2746 4590 2748
rect 4646 2746 4670 2748
rect 4726 2746 4732 2748
rect 4486 2694 4488 2746
rect 4668 2694 4670 2746
rect 4424 2692 4430 2694
rect 4486 2692 4510 2694
rect 4566 2692 4590 2694
rect 4646 2692 4670 2694
rect 4726 2692 4732 2694
rect 4424 2683 4732 2692
rect 5276 2650 5304 5170
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5828 3058 5856 4014
rect 6104 3738 6132 6886
rect 6288 5710 6316 8298
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6380 4690 6408 6734
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6564 5778 6592 6598
rect 6656 6390 6684 8298
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6748 6730 6776 6802
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6644 6384 6696 6390
rect 6644 6326 6696 6332
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6656 4690 6684 4966
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6380 4146 6408 4626
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 6380 3466 6408 4082
rect 7484 3670 7512 5646
rect 7576 5114 7604 8978
rect 7668 8906 7696 13126
rect 7898 13084 8206 13093
rect 7898 13082 7904 13084
rect 7960 13082 7984 13084
rect 8040 13082 8064 13084
rect 8120 13082 8144 13084
rect 8200 13082 8206 13084
rect 7960 13030 7962 13082
rect 8142 13030 8144 13082
rect 7898 13028 7904 13030
rect 7960 13028 7984 13030
rect 8040 13028 8064 13030
rect 8120 13028 8144 13030
rect 8200 13028 8206 13030
rect 7898 13019 8206 13028
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7760 9518 7788 12582
rect 7898 11996 8206 12005
rect 7898 11994 7904 11996
rect 7960 11994 7984 11996
rect 8040 11994 8064 11996
rect 8120 11994 8144 11996
rect 8200 11994 8206 11996
rect 7960 11942 7962 11994
rect 8142 11942 8144 11994
rect 7898 11940 7904 11942
rect 7960 11940 7984 11942
rect 8040 11940 8064 11942
rect 8120 11940 8144 11942
rect 8200 11940 8206 11942
rect 7898 11931 8206 11940
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 7898 10908 8206 10917
rect 7898 10906 7904 10908
rect 7960 10906 7984 10908
rect 8040 10906 8064 10908
rect 8120 10906 8144 10908
rect 8200 10906 8206 10908
rect 7960 10854 7962 10906
rect 8142 10854 8144 10906
rect 7898 10852 7904 10854
rect 7960 10852 7984 10854
rect 8040 10852 8064 10854
rect 8120 10852 8144 10854
rect 8200 10852 8206 10854
rect 7898 10843 8206 10852
rect 7898 9820 8206 9829
rect 7898 9818 7904 9820
rect 7960 9818 7984 9820
rect 8040 9818 8064 9820
rect 8120 9818 8144 9820
rect 8200 9818 8206 9820
rect 7960 9766 7962 9818
rect 8142 9766 8144 9818
rect 7898 9764 7904 9766
rect 7960 9764 7984 9766
rect 8040 9764 8064 9766
rect 8120 9764 8144 9766
rect 8200 9764 8206 9766
rect 7898 9755 8206 9764
rect 8496 9586 8524 11494
rect 9048 10810 9076 14554
rect 9140 13938 9168 15438
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 9324 13870 9352 15438
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9416 13326 9444 13738
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 9508 10742 9536 14350
rect 9600 14074 9628 16390
rect 11372 15804 11680 15813
rect 11372 15802 11378 15804
rect 11434 15802 11458 15804
rect 11514 15802 11538 15804
rect 11594 15802 11618 15804
rect 11674 15802 11680 15804
rect 11434 15750 11436 15802
rect 11616 15750 11618 15802
rect 11372 15748 11378 15750
rect 11434 15748 11458 15750
rect 11514 15748 11538 15750
rect 11594 15748 11618 15750
rect 11674 15748 11680 15750
rect 11372 15739 11680 15748
rect 11716 15706 11744 16390
rect 11808 15910 11836 16510
rect 12452 16114 12480 16526
rect 14846 16348 15154 16357
rect 14846 16346 14852 16348
rect 14908 16346 14932 16348
rect 14988 16346 15012 16348
rect 15068 16346 15092 16348
rect 15148 16346 15154 16348
rect 14908 16294 14910 16346
rect 15090 16294 15092 16346
rect 14846 16292 14852 16294
rect 14908 16292 14932 16294
rect 14988 16292 15012 16294
rect 15068 16292 15092 16294
rect 15148 16292 15154 16294
rect 14846 16283 15154 16292
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 9876 14346 9904 15574
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 10876 14544 10928 14550
rect 10876 14486 10928 14492
rect 10888 14414 10916 14486
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 9864 14340 9916 14346
rect 9864 14282 9916 14288
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9692 14006 9720 14214
rect 9680 14000 9732 14006
rect 9876 13988 9904 14282
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 9876 13960 9996 13988
rect 9680 13942 9732 13948
rect 9692 13326 9720 13942
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9784 13530 9812 13874
rect 9968 13870 9996 13960
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9784 12850 9812 13330
rect 9876 13258 9904 13806
rect 9968 13462 9996 13806
rect 10060 13734 10088 14214
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 10888 13462 10916 14350
rect 11060 14340 11112 14346
rect 11060 14282 11112 14288
rect 11072 13734 11100 14282
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 10876 13456 10928 13462
rect 10876 13398 10928 13404
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 11082 9720 12582
rect 9876 11898 9904 13194
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 10336 10470 10364 11086
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 10062 10364 10406
rect 10612 10130 10640 11494
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10336 9586 10364 9998
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 7656 8900 7708 8906
rect 7656 8842 7708 8848
rect 7898 8732 8206 8741
rect 7898 8730 7904 8732
rect 7960 8730 7984 8732
rect 8040 8730 8064 8732
rect 8120 8730 8144 8732
rect 8200 8730 8206 8732
rect 7960 8678 7962 8730
rect 8142 8678 8144 8730
rect 7898 8676 7904 8678
rect 7960 8676 7984 8678
rect 8040 8676 8064 8678
rect 8120 8676 8144 8678
rect 8200 8676 8206 8678
rect 7898 8667 8206 8676
rect 8496 8498 8524 9522
rect 10704 9518 10732 13126
rect 10796 10742 10824 13126
rect 10888 12850 10916 13398
rect 11072 13394 11100 13670
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 11164 13297 11192 15438
rect 11716 15026 11744 15642
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11372 14716 11680 14725
rect 11372 14714 11378 14716
rect 11434 14714 11458 14716
rect 11514 14714 11538 14716
rect 11594 14714 11618 14716
rect 11674 14714 11680 14716
rect 11434 14662 11436 14714
rect 11616 14662 11618 14714
rect 11372 14660 11378 14662
rect 11434 14660 11458 14662
rect 11514 14660 11538 14662
rect 11594 14660 11618 14662
rect 11674 14660 11680 14662
rect 11372 14651 11680 14660
rect 11808 14618 11836 15846
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11440 14006 11468 14350
rect 11428 14000 11480 14006
rect 11256 13960 11428 13988
rect 11256 13326 11284 13960
rect 11428 13942 11480 13948
rect 11532 13870 11560 14418
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11900 13802 11928 15302
rect 12176 14958 12204 15846
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12348 14340 12400 14346
rect 12348 14282 12400 14288
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 11888 13796 11940 13802
rect 11888 13738 11940 13744
rect 11372 13628 11680 13637
rect 11372 13626 11378 13628
rect 11434 13626 11458 13628
rect 11514 13626 11538 13628
rect 11594 13626 11618 13628
rect 11674 13626 11680 13628
rect 11434 13574 11436 13626
rect 11616 13574 11618 13626
rect 11372 13572 11378 13574
rect 11434 13572 11458 13574
rect 11514 13572 11538 13574
rect 11594 13572 11618 13574
rect 11674 13572 11680 13574
rect 11372 13563 11680 13572
rect 12268 13376 12296 14214
rect 12360 13938 12388 14282
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12348 13388 12400 13394
rect 12268 13348 12348 13376
rect 12348 13330 12400 13336
rect 11244 13320 11296 13326
rect 11150 13288 11206 13297
rect 11244 13262 11296 13268
rect 11150 13223 11206 13232
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11992 12850 12020 13126
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11372 12540 11680 12549
rect 11372 12538 11378 12540
rect 11434 12538 11458 12540
rect 11514 12538 11538 12540
rect 11594 12538 11618 12540
rect 11674 12538 11680 12540
rect 11434 12486 11436 12538
rect 11616 12486 11618 12538
rect 11372 12484 11378 12486
rect 11434 12484 11458 12486
rect 11514 12484 11538 12486
rect 11594 12484 11618 12486
rect 11674 12484 11680 12486
rect 11372 12475 11680 12484
rect 11808 11694 11836 12582
rect 12360 12306 12388 13330
rect 12544 13190 12572 14350
rect 12820 13326 12848 15302
rect 13004 14074 13032 16050
rect 14280 15632 14332 15638
rect 14280 15574 14332 15580
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13188 15162 13216 15302
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13280 14550 13308 15302
rect 13268 14544 13320 14550
rect 13268 14486 13320 14492
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 13280 13734 13308 14486
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12544 12238 12572 13126
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11372 11452 11680 11461
rect 11372 11450 11378 11452
rect 11434 11450 11458 11452
rect 11514 11450 11538 11452
rect 11594 11450 11618 11452
rect 11674 11450 11680 11452
rect 11434 11398 11436 11450
rect 11616 11398 11618 11450
rect 11372 11396 11378 11398
rect 11434 11396 11458 11398
rect 11514 11396 11538 11398
rect 11594 11396 11618 11398
rect 11674 11396 11680 11398
rect 11372 11387 11680 11396
rect 10784 10736 10836 10742
rect 10784 10678 10836 10684
rect 11372 10364 11680 10373
rect 11372 10362 11378 10364
rect 11434 10362 11458 10364
rect 11514 10362 11538 10364
rect 11594 10362 11618 10364
rect 11674 10362 11680 10364
rect 11434 10310 11436 10362
rect 11616 10310 11618 10362
rect 11372 10308 11378 10310
rect 11434 10308 11458 10310
rect 11514 10308 11538 10310
rect 11594 10308 11618 10310
rect 11674 10308 11680 10310
rect 11372 10299 11680 10308
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11164 9654 11192 10066
rect 11716 9654 11744 11494
rect 13280 10810 13308 12174
rect 13648 11354 13676 12718
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13740 10742 13768 13874
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13832 13530 13860 13806
rect 14096 13796 14148 13802
rect 14096 13738 14148 13744
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13924 11218 13952 12582
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 14108 11150 14136 13738
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14200 12850 14228 13194
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 13728 10736 13780 10742
rect 13728 10678 13780 10684
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 12716 9988 12768 9994
rect 12716 9930 12768 9936
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 11372 9276 11680 9285
rect 11372 9274 11378 9276
rect 11434 9274 11458 9276
rect 11514 9274 11538 9276
rect 11594 9274 11618 9276
rect 11674 9274 11680 9276
rect 11434 9222 11436 9274
rect 11616 9222 11618 9274
rect 11372 9220 11378 9222
rect 11434 9220 11458 9222
rect 11514 9220 11538 9222
rect 11594 9220 11618 9222
rect 11674 9220 11680 9222
rect 11372 9211 11680 9220
rect 12728 9178 12756 9930
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13740 9654 13768 9862
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 14016 9382 14044 10202
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8496 7954 8524 8434
rect 9784 8090 9812 8502
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7668 7206 7696 7754
rect 7898 7644 8206 7653
rect 7898 7642 7904 7644
rect 7960 7642 7984 7644
rect 8040 7642 8064 7644
rect 8120 7642 8144 7644
rect 8200 7642 8206 7644
rect 7960 7590 7962 7642
rect 8142 7590 8144 7642
rect 7898 7588 7904 7590
rect 7960 7588 7984 7590
rect 8040 7588 8064 7590
rect 8120 7588 8144 7590
rect 8200 7588 8206 7590
rect 7898 7579 8206 7588
rect 8496 7410 8524 7890
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 10060 7342 10088 8910
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11256 7954 11284 8230
rect 11372 8188 11680 8197
rect 11372 8186 11378 8188
rect 11434 8186 11458 8188
rect 11514 8186 11538 8188
rect 11594 8186 11618 8188
rect 11674 8186 11680 8188
rect 11434 8134 11436 8186
rect 11616 8134 11618 8186
rect 11372 8132 11378 8134
rect 11434 8132 11458 8134
rect 11514 8132 11538 8134
rect 11594 8132 11618 8134
rect 11674 8132 11680 8134
rect 11372 8123 11680 8132
rect 12360 8090 12388 8502
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11348 7546 11376 7890
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12268 7546 12296 7754
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 14016 7478 14044 8366
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 14108 8090 14136 8298
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14004 7472 14056 7478
rect 14004 7414 14056 7420
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 10784 7268 10836 7274
rect 10784 7210 10836 7216
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7668 5302 7696 7142
rect 10796 6866 10824 7210
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 11372 7100 11680 7109
rect 11372 7098 11378 7100
rect 11434 7098 11458 7100
rect 11514 7098 11538 7100
rect 11594 7098 11618 7100
rect 11674 7098 11680 7100
rect 11434 7046 11436 7098
rect 11616 7046 11618 7098
rect 11372 7044 11378 7046
rect 11434 7044 11458 7046
rect 11514 7044 11538 7046
rect 11594 7044 11618 7046
rect 11674 7044 11680 7046
rect 11372 7035 11680 7044
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 10324 6792 10376 6798
rect 7746 6760 7802 6769
rect 10324 6734 10376 6740
rect 7746 6695 7802 6704
rect 7760 6322 7788 6695
rect 7898 6556 8206 6565
rect 7898 6554 7904 6556
rect 7960 6554 7984 6556
rect 8040 6554 8064 6556
rect 8120 6554 8144 6556
rect 8200 6554 8206 6556
rect 7960 6502 7962 6554
rect 8142 6502 8144 6554
rect 7898 6500 7904 6502
rect 7960 6500 7984 6502
rect 8040 6500 8064 6502
rect 8120 6500 8144 6502
rect 8200 6500 8206 6502
rect 7898 6491 8206 6500
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8588 5778 8616 6190
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8680 5914 8708 6054
rect 8956 5914 8984 6190
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 10336 5778 10364 6734
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 10704 5778 10732 6666
rect 11164 6322 11192 6666
rect 11256 6458 11284 6802
rect 13188 6730 13216 7142
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14108 6905 14136 6938
rect 14094 6896 14150 6905
rect 14094 6831 14150 6840
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 14096 6724 14148 6730
rect 14096 6666 14148 6672
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 12820 6390 12848 6598
rect 12808 6384 12860 6390
rect 12808 6326 12860 6332
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 11072 5846 11100 6258
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 11372 6012 11680 6021
rect 11372 6010 11378 6012
rect 11434 6010 11458 6012
rect 11514 6010 11538 6012
rect 11594 6010 11618 6012
rect 11674 6010 11680 6012
rect 11434 5958 11436 6010
rect 11616 5958 11618 6010
rect 11372 5956 11378 5958
rect 11434 5956 11458 5958
rect 11514 5956 11538 5958
rect 11594 5956 11618 5958
rect 11674 5956 11680 5958
rect 11372 5947 11680 5956
rect 12820 5914 12848 6054
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 7898 5468 8206 5477
rect 7898 5466 7904 5468
rect 7960 5466 7984 5468
rect 8040 5466 8064 5468
rect 8120 5466 8144 5468
rect 8200 5466 8206 5468
rect 7960 5414 7962 5466
rect 8142 5414 8144 5466
rect 7898 5412 7904 5414
rect 7960 5412 7984 5414
rect 8040 5412 8064 5414
rect 8120 5412 8144 5414
rect 8200 5412 8206 5414
rect 7898 5403 8206 5412
rect 8588 5370 8616 5714
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 9968 5234 9996 5578
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 8116 5160 8168 5166
rect 7576 5086 7696 5114
rect 8116 5102 8168 5108
rect 7668 4554 7696 5086
rect 8128 4826 8156 5102
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 10336 4690 10364 5714
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11372 4924 11680 4933
rect 11372 4922 11378 4924
rect 11434 4922 11458 4924
rect 11514 4922 11538 4924
rect 11594 4922 11618 4924
rect 11674 4922 11680 4924
rect 11434 4870 11436 4922
rect 11616 4870 11618 4922
rect 11372 4868 11378 4870
rect 11434 4868 11458 4870
rect 11514 4868 11538 4870
rect 11594 4868 11618 4870
rect 11674 4868 11680 4870
rect 11372 4859 11680 4868
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 7898 4380 8206 4389
rect 7898 4378 7904 4380
rect 7960 4378 7984 4380
rect 8040 4378 8064 4380
rect 8120 4378 8144 4380
rect 8200 4378 8206 4380
rect 7960 4326 7962 4378
rect 8142 4326 8144 4378
rect 7898 4324 7904 4326
rect 7960 4324 7984 4326
rect 8040 4324 8064 4326
rect 8120 4324 8144 4326
rect 8200 4324 8206 4326
rect 7898 4315 8206 4324
rect 10336 4146 10364 4626
rect 10600 4548 10652 4554
rect 10600 4490 10652 4496
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 6564 3058 6592 3402
rect 8036 3398 8064 3878
rect 10336 3602 10364 4082
rect 10612 4078 10640 4490
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 7760 2990 7788 3334
rect 7898 3292 8206 3301
rect 7898 3290 7904 3292
rect 7960 3290 7984 3292
rect 8040 3290 8064 3292
rect 8120 3290 8144 3292
rect 8200 3290 8206 3292
rect 7960 3238 7962 3290
rect 8142 3238 8144 3290
rect 7898 3236 7904 3238
rect 7960 3236 7984 3238
rect 8040 3236 8064 3238
rect 8120 3236 8144 3238
rect 8200 3236 8206 3238
rect 7898 3227 8206 3236
rect 8496 3126 8524 3470
rect 10336 3194 10364 3538
rect 10600 3460 10652 3466
rect 10600 3402 10652 3408
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 10612 3194 10640 3402
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 8484 3120 8536 3126
rect 8484 3062 8536 3068
rect 10796 3058 10824 3402
rect 10980 3126 11008 4626
rect 11716 4214 11744 4966
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 12912 3942 12940 6190
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 13096 4826 13124 5578
rect 13188 5098 13216 6258
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13176 5092 13228 5098
rect 13176 5034 13228 5040
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 13556 4622 13584 5510
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13556 4486 13584 4558
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13740 4214 13768 4966
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 11372 3836 11680 3845
rect 11372 3834 11378 3836
rect 11434 3834 11458 3836
rect 11514 3834 11538 3836
rect 11594 3834 11618 3836
rect 11674 3834 11680 3836
rect 11434 3782 11436 3834
rect 11616 3782 11618 3834
rect 11372 3780 11378 3782
rect 11434 3780 11458 3782
rect 11514 3780 11538 3782
rect 11594 3780 11618 3782
rect 11674 3780 11680 3782
rect 11372 3771 11680 3780
rect 14016 3670 14044 6258
rect 14108 5166 14136 6666
rect 14200 6458 14228 12786
rect 14292 9518 14320 15574
rect 14846 15260 15154 15269
rect 14846 15258 14852 15260
rect 14908 15258 14932 15260
rect 14988 15258 15012 15260
rect 15068 15258 15092 15260
rect 15148 15258 15154 15260
rect 14908 15206 14910 15258
rect 15090 15206 15092 15258
rect 14846 15204 14852 15206
rect 14908 15204 14932 15206
rect 14988 15204 15012 15206
rect 15068 15204 15092 15206
rect 15148 15204 15154 15206
rect 14846 15195 15154 15204
rect 14846 14172 15154 14181
rect 14846 14170 14852 14172
rect 14908 14170 14932 14172
rect 14988 14170 15012 14172
rect 15068 14170 15092 14172
rect 15148 14170 15154 14172
rect 14908 14118 14910 14170
rect 15090 14118 15092 14170
rect 14846 14116 14852 14118
rect 14908 14116 14932 14118
rect 14988 14116 15012 14118
rect 15068 14116 15092 14118
rect 15148 14116 15154 14118
rect 14846 14107 15154 14116
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 14384 12986 14412 13262
rect 14846 13084 15154 13093
rect 14846 13082 14852 13084
rect 14908 13082 14932 13084
rect 14988 13082 15012 13084
rect 15068 13082 15092 13084
rect 15148 13082 15154 13084
rect 14908 13030 14910 13082
rect 15090 13030 15092 13082
rect 14846 13028 14852 13030
rect 14908 13028 14932 13030
rect 14988 13028 15012 13030
rect 15068 13028 15092 13030
rect 15148 13028 15154 13030
rect 14846 13019 15154 13028
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14660 10062 14688 11086
rect 14752 10674 14780 12038
rect 14846 11996 15154 12005
rect 14846 11994 14852 11996
rect 14908 11994 14932 11996
rect 14988 11994 15012 11996
rect 15068 11994 15092 11996
rect 15148 11994 15154 11996
rect 14908 11942 14910 11994
rect 15090 11942 15092 11994
rect 14846 11940 14852 11942
rect 14908 11940 14932 11942
rect 14988 11940 15012 11942
rect 15068 11940 15092 11942
rect 15148 11940 15154 11942
rect 14846 11931 15154 11940
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14844 11354 14872 11698
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14846 10908 15154 10917
rect 14846 10906 14852 10908
rect 14908 10906 14932 10908
rect 14988 10906 15012 10908
rect 15068 10906 15092 10908
rect 15148 10906 15154 10908
rect 14908 10854 14910 10906
rect 15090 10854 15092 10906
rect 14846 10852 14852 10854
rect 14908 10852 14932 10854
rect 14988 10852 15012 10854
rect 15068 10852 15092 10854
rect 15148 10852 15154 10854
rect 14846 10843 15154 10852
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14846 9820 15154 9829
rect 14846 9818 14852 9820
rect 14908 9818 14932 9820
rect 14988 9818 15012 9820
rect 15068 9818 15092 9820
rect 15148 9818 15154 9820
rect 14908 9766 14910 9818
rect 15090 9766 15092 9818
rect 14846 9764 14852 9766
rect 14908 9764 14932 9766
rect 14988 9764 15012 9766
rect 15068 9764 15092 9766
rect 15148 9764 15154 9766
rect 14846 9755 15154 9764
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14292 5386 14320 7822
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14200 5358 14320 5386
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 14200 4826 14228 5358
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14292 4622 14320 5170
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14384 4078 14412 6734
rect 14476 6390 14504 7822
rect 14660 7342 14688 9590
rect 15304 9586 15332 13262
rect 15580 12714 15608 13466
rect 15568 12708 15620 12714
rect 15568 12650 15620 12656
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14752 8498 14780 8910
rect 14846 8732 15154 8741
rect 14846 8730 14852 8732
rect 14908 8730 14932 8732
rect 14988 8730 15012 8732
rect 15068 8730 15092 8732
rect 15148 8730 15154 8732
rect 14908 8678 14910 8730
rect 15090 8678 15092 8730
rect 14846 8676 14852 8678
rect 14908 8676 14932 8678
rect 14988 8676 15012 8678
rect 15068 8676 15092 8678
rect 15148 8676 15154 8678
rect 14846 8667 15154 8676
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14752 7818 14780 8434
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 14752 7410 14780 7754
rect 14846 7644 15154 7653
rect 14846 7642 14852 7644
rect 14908 7642 14932 7644
rect 14988 7642 15012 7644
rect 15068 7642 15092 7644
rect 15148 7642 15154 7644
rect 14908 7590 14910 7642
rect 15090 7590 15092 7642
rect 14846 7588 14852 7590
rect 14908 7588 14932 7590
rect 14988 7588 15012 7590
rect 15068 7588 15092 7590
rect 15148 7588 15154 7590
rect 14846 7579 15154 7588
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14464 6384 14516 6390
rect 14464 6326 14516 6332
rect 14568 6118 14596 6598
rect 14660 6458 14688 7278
rect 15304 6914 15332 9522
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15396 7886 15424 9318
rect 15580 8090 15608 12650
rect 18156 12442 18184 27270
rect 21794 27228 22102 27237
rect 21794 27226 21800 27228
rect 21856 27226 21880 27228
rect 21936 27226 21960 27228
rect 22016 27226 22040 27228
rect 22096 27226 22102 27228
rect 21856 27174 21858 27226
rect 22038 27174 22040 27226
rect 21794 27172 21800 27174
rect 21856 27172 21880 27174
rect 21936 27172 21960 27174
rect 22016 27172 22040 27174
rect 22096 27172 22102 27174
rect 21794 27163 22102 27172
rect 18320 26684 18628 26693
rect 18320 26682 18326 26684
rect 18382 26682 18406 26684
rect 18462 26682 18486 26684
rect 18542 26682 18566 26684
rect 18622 26682 18628 26684
rect 18382 26630 18384 26682
rect 18564 26630 18566 26682
rect 18320 26628 18326 26630
rect 18382 26628 18406 26630
rect 18462 26628 18486 26630
rect 18542 26628 18566 26630
rect 18622 26628 18628 26630
rect 18320 26619 18628 26628
rect 25268 26684 25576 26693
rect 25268 26682 25274 26684
rect 25330 26682 25354 26684
rect 25410 26682 25434 26684
rect 25490 26682 25514 26684
rect 25570 26682 25576 26684
rect 25330 26630 25332 26682
rect 25512 26630 25514 26682
rect 25268 26628 25274 26630
rect 25330 26628 25354 26630
rect 25410 26628 25434 26630
rect 25490 26628 25514 26630
rect 25570 26628 25576 26630
rect 25268 26619 25576 26628
rect 21794 26140 22102 26149
rect 21794 26138 21800 26140
rect 21856 26138 21880 26140
rect 21936 26138 21960 26140
rect 22016 26138 22040 26140
rect 22096 26138 22102 26140
rect 21856 26086 21858 26138
rect 22038 26086 22040 26138
rect 21794 26084 21800 26086
rect 21856 26084 21880 26086
rect 21936 26084 21960 26086
rect 22016 26084 22040 26086
rect 22096 26084 22102 26086
rect 21794 26075 22102 26084
rect 18320 25596 18628 25605
rect 18320 25594 18326 25596
rect 18382 25594 18406 25596
rect 18462 25594 18486 25596
rect 18542 25594 18566 25596
rect 18622 25594 18628 25596
rect 18382 25542 18384 25594
rect 18564 25542 18566 25594
rect 18320 25540 18326 25542
rect 18382 25540 18406 25542
rect 18462 25540 18486 25542
rect 18542 25540 18566 25542
rect 18622 25540 18628 25542
rect 18320 25531 18628 25540
rect 25268 25596 25576 25605
rect 25268 25594 25274 25596
rect 25330 25594 25354 25596
rect 25410 25594 25434 25596
rect 25490 25594 25514 25596
rect 25570 25594 25576 25596
rect 25330 25542 25332 25594
rect 25512 25542 25514 25594
rect 25268 25540 25274 25542
rect 25330 25540 25354 25542
rect 25410 25540 25434 25542
rect 25490 25540 25514 25542
rect 25570 25540 25576 25542
rect 25268 25531 25576 25540
rect 21794 25052 22102 25061
rect 21794 25050 21800 25052
rect 21856 25050 21880 25052
rect 21936 25050 21960 25052
rect 22016 25050 22040 25052
rect 22096 25050 22102 25052
rect 21856 24998 21858 25050
rect 22038 24998 22040 25050
rect 21794 24996 21800 24998
rect 21856 24996 21880 24998
rect 21936 24996 21960 24998
rect 22016 24996 22040 24998
rect 22096 24996 22102 24998
rect 21794 24987 22102 24996
rect 18320 24508 18628 24517
rect 18320 24506 18326 24508
rect 18382 24506 18406 24508
rect 18462 24506 18486 24508
rect 18542 24506 18566 24508
rect 18622 24506 18628 24508
rect 18382 24454 18384 24506
rect 18564 24454 18566 24506
rect 18320 24452 18326 24454
rect 18382 24452 18406 24454
rect 18462 24452 18486 24454
rect 18542 24452 18566 24454
rect 18622 24452 18628 24454
rect 18320 24443 18628 24452
rect 25268 24508 25576 24517
rect 25268 24506 25274 24508
rect 25330 24506 25354 24508
rect 25410 24506 25434 24508
rect 25490 24506 25514 24508
rect 25570 24506 25576 24508
rect 25330 24454 25332 24506
rect 25512 24454 25514 24506
rect 25268 24452 25274 24454
rect 25330 24452 25354 24454
rect 25410 24452 25434 24454
rect 25490 24452 25514 24454
rect 25570 24452 25576 24454
rect 25268 24443 25576 24452
rect 21794 23964 22102 23973
rect 21794 23962 21800 23964
rect 21856 23962 21880 23964
rect 21936 23962 21960 23964
rect 22016 23962 22040 23964
rect 22096 23962 22102 23964
rect 21856 23910 21858 23962
rect 22038 23910 22040 23962
rect 21794 23908 21800 23910
rect 21856 23908 21880 23910
rect 21936 23908 21960 23910
rect 22016 23908 22040 23910
rect 22096 23908 22102 23910
rect 21794 23899 22102 23908
rect 18320 23420 18628 23429
rect 18320 23418 18326 23420
rect 18382 23418 18406 23420
rect 18462 23418 18486 23420
rect 18542 23418 18566 23420
rect 18622 23418 18628 23420
rect 18382 23366 18384 23418
rect 18564 23366 18566 23418
rect 18320 23364 18326 23366
rect 18382 23364 18406 23366
rect 18462 23364 18486 23366
rect 18542 23364 18566 23366
rect 18622 23364 18628 23366
rect 18320 23355 18628 23364
rect 25268 23420 25576 23429
rect 25268 23418 25274 23420
rect 25330 23418 25354 23420
rect 25410 23418 25434 23420
rect 25490 23418 25514 23420
rect 25570 23418 25576 23420
rect 25330 23366 25332 23418
rect 25512 23366 25514 23418
rect 25268 23364 25274 23366
rect 25330 23364 25354 23366
rect 25410 23364 25434 23366
rect 25490 23364 25514 23366
rect 25570 23364 25576 23366
rect 25268 23355 25576 23364
rect 21794 22876 22102 22885
rect 21794 22874 21800 22876
rect 21856 22874 21880 22876
rect 21936 22874 21960 22876
rect 22016 22874 22040 22876
rect 22096 22874 22102 22876
rect 21856 22822 21858 22874
rect 22038 22822 22040 22874
rect 21794 22820 21800 22822
rect 21856 22820 21880 22822
rect 21936 22820 21960 22822
rect 22016 22820 22040 22822
rect 22096 22820 22102 22822
rect 21794 22811 22102 22820
rect 18320 22332 18628 22341
rect 18320 22330 18326 22332
rect 18382 22330 18406 22332
rect 18462 22330 18486 22332
rect 18542 22330 18566 22332
rect 18622 22330 18628 22332
rect 18382 22278 18384 22330
rect 18564 22278 18566 22330
rect 18320 22276 18326 22278
rect 18382 22276 18406 22278
rect 18462 22276 18486 22278
rect 18542 22276 18566 22278
rect 18622 22276 18628 22278
rect 18320 22267 18628 22276
rect 25268 22332 25576 22341
rect 25268 22330 25274 22332
rect 25330 22330 25354 22332
rect 25410 22330 25434 22332
rect 25490 22330 25514 22332
rect 25570 22330 25576 22332
rect 25330 22278 25332 22330
rect 25512 22278 25514 22330
rect 25268 22276 25274 22278
rect 25330 22276 25354 22278
rect 25410 22276 25434 22278
rect 25490 22276 25514 22278
rect 25570 22276 25576 22278
rect 25268 22267 25576 22276
rect 21794 21788 22102 21797
rect 21794 21786 21800 21788
rect 21856 21786 21880 21788
rect 21936 21786 21960 21788
rect 22016 21786 22040 21788
rect 22096 21786 22102 21788
rect 21856 21734 21858 21786
rect 22038 21734 22040 21786
rect 21794 21732 21800 21734
rect 21856 21732 21880 21734
rect 21936 21732 21960 21734
rect 22016 21732 22040 21734
rect 22096 21732 22102 21734
rect 21794 21723 22102 21732
rect 18320 21244 18628 21253
rect 18320 21242 18326 21244
rect 18382 21242 18406 21244
rect 18462 21242 18486 21244
rect 18542 21242 18566 21244
rect 18622 21242 18628 21244
rect 18382 21190 18384 21242
rect 18564 21190 18566 21242
rect 18320 21188 18326 21190
rect 18382 21188 18406 21190
rect 18462 21188 18486 21190
rect 18542 21188 18566 21190
rect 18622 21188 18628 21190
rect 18320 21179 18628 21188
rect 25268 21244 25576 21253
rect 25268 21242 25274 21244
rect 25330 21242 25354 21244
rect 25410 21242 25434 21244
rect 25490 21242 25514 21244
rect 25570 21242 25576 21244
rect 25330 21190 25332 21242
rect 25512 21190 25514 21242
rect 25268 21188 25274 21190
rect 25330 21188 25354 21190
rect 25410 21188 25434 21190
rect 25490 21188 25514 21190
rect 25570 21188 25576 21190
rect 25268 21179 25576 21188
rect 21794 20700 22102 20709
rect 21794 20698 21800 20700
rect 21856 20698 21880 20700
rect 21936 20698 21960 20700
rect 22016 20698 22040 20700
rect 22096 20698 22102 20700
rect 21856 20646 21858 20698
rect 22038 20646 22040 20698
rect 21794 20644 21800 20646
rect 21856 20644 21880 20646
rect 21936 20644 21960 20646
rect 22016 20644 22040 20646
rect 22096 20644 22102 20646
rect 21794 20635 22102 20644
rect 18320 20156 18628 20165
rect 18320 20154 18326 20156
rect 18382 20154 18406 20156
rect 18462 20154 18486 20156
rect 18542 20154 18566 20156
rect 18622 20154 18628 20156
rect 18382 20102 18384 20154
rect 18564 20102 18566 20154
rect 18320 20100 18326 20102
rect 18382 20100 18406 20102
rect 18462 20100 18486 20102
rect 18542 20100 18566 20102
rect 18622 20100 18628 20102
rect 18320 20091 18628 20100
rect 25268 20156 25576 20165
rect 25268 20154 25274 20156
rect 25330 20154 25354 20156
rect 25410 20154 25434 20156
rect 25490 20154 25514 20156
rect 25570 20154 25576 20156
rect 25330 20102 25332 20154
rect 25512 20102 25514 20154
rect 25268 20100 25274 20102
rect 25330 20100 25354 20102
rect 25410 20100 25434 20102
rect 25490 20100 25514 20102
rect 25570 20100 25576 20102
rect 25268 20091 25576 20100
rect 21794 19612 22102 19621
rect 21794 19610 21800 19612
rect 21856 19610 21880 19612
rect 21936 19610 21960 19612
rect 22016 19610 22040 19612
rect 22096 19610 22102 19612
rect 21856 19558 21858 19610
rect 22038 19558 22040 19610
rect 21794 19556 21800 19558
rect 21856 19556 21880 19558
rect 21936 19556 21960 19558
rect 22016 19556 22040 19558
rect 22096 19556 22102 19558
rect 21794 19547 22102 19556
rect 18320 19068 18628 19077
rect 18320 19066 18326 19068
rect 18382 19066 18406 19068
rect 18462 19066 18486 19068
rect 18542 19066 18566 19068
rect 18622 19066 18628 19068
rect 18382 19014 18384 19066
rect 18564 19014 18566 19066
rect 18320 19012 18326 19014
rect 18382 19012 18406 19014
rect 18462 19012 18486 19014
rect 18542 19012 18566 19014
rect 18622 19012 18628 19014
rect 18320 19003 18628 19012
rect 25268 19068 25576 19077
rect 25268 19066 25274 19068
rect 25330 19066 25354 19068
rect 25410 19066 25434 19068
rect 25490 19066 25514 19068
rect 25570 19066 25576 19068
rect 25330 19014 25332 19066
rect 25512 19014 25514 19066
rect 25268 19012 25274 19014
rect 25330 19012 25354 19014
rect 25410 19012 25434 19014
rect 25490 19012 25514 19014
rect 25570 19012 25576 19014
rect 25268 19003 25576 19012
rect 21794 18524 22102 18533
rect 21794 18522 21800 18524
rect 21856 18522 21880 18524
rect 21936 18522 21960 18524
rect 22016 18522 22040 18524
rect 22096 18522 22102 18524
rect 21856 18470 21858 18522
rect 22038 18470 22040 18522
rect 21794 18468 21800 18470
rect 21856 18468 21880 18470
rect 21936 18468 21960 18470
rect 22016 18468 22040 18470
rect 22096 18468 22102 18470
rect 21794 18459 22102 18468
rect 18320 17980 18628 17989
rect 18320 17978 18326 17980
rect 18382 17978 18406 17980
rect 18462 17978 18486 17980
rect 18542 17978 18566 17980
rect 18622 17978 18628 17980
rect 18382 17926 18384 17978
rect 18564 17926 18566 17978
rect 18320 17924 18326 17926
rect 18382 17924 18406 17926
rect 18462 17924 18486 17926
rect 18542 17924 18566 17926
rect 18622 17924 18628 17926
rect 18320 17915 18628 17924
rect 25268 17980 25576 17989
rect 25268 17978 25274 17980
rect 25330 17978 25354 17980
rect 25410 17978 25434 17980
rect 25490 17978 25514 17980
rect 25570 17978 25576 17980
rect 25330 17926 25332 17978
rect 25512 17926 25514 17978
rect 25268 17924 25274 17926
rect 25330 17924 25354 17926
rect 25410 17924 25434 17926
rect 25490 17924 25514 17926
rect 25570 17924 25576 17926
rect 25268 17915 25576 17924
rect 21794 17436 22102 17445
rect 21794 17434 21800 17436
rect 21856 17434 21880 17436
rect 21936 17434 21960 17436
rect 22016 17434 22040 17436
rect 22096 17434 22102 17436
rect 21856 17382 21858 17434
rect 22038 17382 22040 17434
rect 21794 17380 21800 17382
rect 21856 17380 21880 17382
rect 21936 17380 21960 17382
rect 22016 17380 22040 17382
rect 22096 17380 22102 17382
rect 21794 17371 22102 17380
rect 28172 17196 28224 17202
rect 28172 17138 28224 17144
rect 28184 17105 28212 17138
rect 28170 17096 28226 17105
rect 28170 17031 28226 17040
rect 27988 16992 28040 16998
rect 27988 16934 28040 16940
rect 18320 16892 18628 16901
rect 18320 16890 18326 16892
rect 18382 16890 18406 16892
rect 18462 16890 18486 16892
rect 18542 16890 18566 16892
rect 18622 16890 18628 16892
rect 18382 16838 18384 16890
rect 18564 16838 18566 16890
rect 18320 16836 18326 16838
rect 18382 16836 18406 16838
rect 18462 16836 18486 16838
rect 18542 16836 18566 16838
rect 18622 16836 18628 16838
rect 18320 16827 18628 16836
rect 25268 16892 25576 16901
rect 25268 16890 25274 16892
rect 25330 16890 25354 16892
rect 25410 16890 25434 16892
rect 25490 16890 25514 16892
rect 25570 16890 25576 16892
rect 25330 16838 25332 16890
rect 25512 16838 25514 16890
rect 25268 16836 25274 16838
rect 25330 16836 25354 16838
rect 25410 16836 25434 16838
rect 25490 16836 25514 16838
rect 25570 16836 25576 16838
rect 25268 16827 25576 16836
rect 21794 16348 22102 16357
rect 21794 16346 21800 16348
rect 21856 16346 21880 16348
rect 21936 16346 21960 16348
rect 22016 16346 22040 16348
rect 22096 16346 22102 16348
rect 21856 16294 21858 16346
rect 22038 16294 22040 16346
rect 21794 16292 21800 16294
rect 21856 16292 21880 16294
rect 21936 16292 21960 16294
rect 22016 16292 22040 16294
rect 22096 16292 22102 16294
rect 21794 16283 22102 16292
rect 18320 15804 18628 15813
rect 18320 15802 18326 15804
rect 18382 15802 18406 15804
rect 18462 15802 18486 15804
rect 18542 15802 18566 15804
rect 18622 15802 18628 15804
rect 18382 15750 18384 15802
rect 18564 15750 18566 15802
rect 18320 15748 18326 15750
rect 18382 15748 18406 15750
rect 18462 15748 18486 15750
rect 18542 15748 18566 15750
rect 18622 15748 18628 15750
rect 18320 15739 18628 15748
rect 25268 15804 25576 15813
rect 25268 15802 25274 15804
rect 25330 15802 25354 15804
rect 25410 15802 25434 15804
rect 25490 15802 25514 15804
rect 25570 15802 25576 15804
rect 25330 15750 25332 15802
rect 25512 15750 25514 15802
rect 25268 15748 25274 15750
rect 25330 15748 25354 15750
rect 25410 15748 25434 15750
rect 25490 15748 25514 15750
rect 25570 15748 25576 15750
rect 25268 15739 25576 15748
rect 21794 15260 22102 15269
rect 21794 15258 21800 15260
rect 21856 15258 21880 15260
rect 21936 15258 21960 15260
rect 22016 15258 22040 15260
rect 22096 15258 22102 15260
rect 21856 15206 21858 15258
rect 22038 15206 22040 15258
rect 21794 15204 21800 15206
rect 21856 15204 21880 15206
rect 21936 15204 21960 15206
rect 22016 15204 22040 15206
rect 22096 15204 22102 15206
rect 21794 15195 22102 15204
rect 28000 14822 28028 16934
rect 27988 14816 28040 14822
rect 27988 14758 28040 14764
rect 18320 14716 18628 14725
rect 18320 14714 18326 14716
rect 18382 14714 18406 14716
rect 18462 14714 18486 14716
rect 18542 14714 18566 14716
rect 18622 14714 18628 14716
rect 18382 14662 18384 14714
rect 18564 14662 18566 14714
rect 18320 14660 18326 14662
rect 18382 14660 18406 14662
rect 18462 14660 18486 14662
rect 18542 14660 18566 14662
rect 18622 14660 18628 14662
rect 18320 14651 18628 14660
rect 25268 14716 25576 14725
rect 25268 14714 25274 14716
rect 25330 14714 25354 14716
rect 25410 14714 25434 14716
rect 25490 14714 25514 14716
rect 25570 14714 25576 14716
rect 25330 14662 25332 14714
rect 25512 14662 25514 14714
rect 25268 14660 25274 14662
rect 25330 14660 25354 14662
rect 25410 14660 25434 14662
rect 25490 14660 25514 14662
rect 25570 14660 25576 14662
rect 25268 14651 25576 14660
rect 21794 14172 22102 14181
rect 21794 14170 21800 14172
rect 21856 14170 21880 14172
rect 21936 14170 21960 14172
rect 22016 14170 22040 14172
rect 22096 14170 22102 14172
rect 21856 14118 21858 14170
rect 22038 14118 22040 14170
rect 21794 14116 21800 14118
rect 21856 14116 21880 14118
rect 21936 14116 21960 14118
rect 22016 14116 22040 14118
rect 22096 14116 22102 14118
rect 21794 14107 22102 14116
rect 18320 13628 18628 13637
rect 18320 13626 18326 13628
rect 18382 13626 18406 13628
rect 18462 13626 18486 13628
rect 18542 13626 18566 13628
rect 18622 13626 18628 13628
rect 18382 13574 18384 13626
rect 18564 13574 18566 13626
rect 18320 13572 18326 13574
rect 18382 13572 18406 13574
rect 18462 13572 18486 13574
rect 18542 13572 18566 13574
rect 18622 13572 18628 13574
rect 18320 13563 18628 13572
rect 25268 13628 25576 13637
rect 25268 13626 25274 13628
rect 25330 13626 25354 13628
rect 25410 13626 25434 13628
rect 25490 13626 25514 13628
rect 25570 13626 25576 13628
rect 25330 13574 25332 13626
rect 25512 13574 25514 13626
rect 25268 13572 25274 13574
rect 25330 13572 25354 13574
rect 25410 13572 25434 13574
rect 25490 13572 25514 13574
rect 25570 13572 25576 13574
rect 25268 13563 25576 13572
rect 21794 13084 22102 13093
rect 21794 13082 21800 13084
rect 21856 13082 21880 13084
rect 21936 13082 21960 13084
rect 22016 13082 22040 13084
rect 22096 13082 22102 13084
rect 21856 13030 21858 13082
rect 22038 13030 22040 13082
rect 21794 13028 21800 13030
rect 21856 13028 21880 13030
rect 21936 13028 21960 13030
rect 22016 13028 22040 13030
rect 22096 13028 22102 13030
rect 21794 13019 22102 13028
rect 18320 12540 18628 12549
rect 18320 12538 18326 12540
rect 18382 12538 18406 12540
rect 18462 12538 18486 12540
rect 18542 12538 18566 12540
rect 18622 12538 18628 12540
rect 18382 12486 18384 12538
rect 18564 12486 18566 12538
rect 18320 12484 18326 12486
rect 18382 12484 18406 12486
rect 18462 12484 18486 12486
rect 18542 12484 18566 12486
rect 18622 12484 18628 12486
rect 18320 12475 18628 12484
rect 25268 12540 25576 12549
rect 25268 12538 25274 12540
rect 25330 12538 25354 12540
rect 25410 12538 25434 12540
rect 25490 12538 25514 12540
rect 25570 12538 25576 12540
rect 25330 12486 25332 12538
rect 25512 12486 25514 12538
rect 25268 12484 25274 12486
rect 25330 12484 25354 12486
rect 25410 12484 25434 12486
rect 25490 12484 25514 12486
rect 25570 12484 25576 12486
rect 25268 12475 25576 12484
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 21794 11996 22102 12005
rect 21794 11994 21800 11996
rect 21856 11994 21880 11996
rect 21936 11994 21960 11996
rect 22016 11994 22040 11996
rect 22096 11994 22102 11996
rect 21856 11942 21858 11994
rect 22038 11942 22040 11994
rect 21794 11940 21800 11942
rect 21856 11940 21880 11942
rect 21936 11940 21960 11942
rect 22016 11940 22040 11942
rect 22096 11940 22102 11942
rect 21794 11931 22102 11940
rect 18320 11452 18628 11461
rect 18320 11450 18326 11452
rect 18382 11450 18406 11452
rect 18462 11450 18486 11452
rect 18542 11450 18566 11452
rect 18622 11450 18628 11452
rect 18382 11398 18384 11450
rect 18564 11398 18566 11450
rect 18320 11396 18326 11398
rect 18382 11396 18406 11398
rect 18462 11396 18486 11398
rect 18542 11396 18566 11398
rect 18622 11396 18628 11398
rect 18320 11387 18628 11396
rect 25268 11452 25576 11461
rect 25268 11450 25274 11452
rect 25330 11450 25354 11452
rect 25410 11450 25434 11452
rect 25490 11450 25514 11452
rect 25570 11450 25576 11452
rect 25330 11398 25332 11450
rect 25512 11398 25514 11450
rect 25268 11396 25274 11398
rect 25330 11396 25354 11398
rect 25410 11396 25434 11398
rect 25490 11396 25514 11398
rect 25570 11396 25576 11398
rect 25268 11387 25576 11396
rect 21794 10908 22102 10917
rect 21794 10906 21800 10908
rect 21856 10906 21880 10908
rect 21936 10906 21960 10908
rect 22016 10906 22040 10908
rect 22096 10906 22102 10908
rect 21856 10854 21858 10906
rect 22038 10854 22040 10906
rect 21794 10852 21800 10854
rect 21856 10852 21880 10854
rect 21936 10852 21960 10854
rect 22016 10852 22040 10854
rect 22096 10852 22102 10854
rect 21794 10843 22102 10852
rect 18320 10364 18628 10373
rect 18320 10362 18326 10364
rect 18382 10362 18406 10364
rect 18462 10362 18486 10364
rect 18542 10362 18566 10364
rect 18622 10362 18628 10364
rect 18382 10310 18384 10362
rect 18564 10310 18566 10362
rect 18320 10308 18326 10310
rect 18382 10308 18406 10310
rect 18462 10308 18486 10310
rect 18542 10308 18566 10310
rect 18622 10308 18628 10310
rect 18320 10299 18628 10308
rect 25268 10364 25576 10373
rect 25268 10362 25274 10364
rect 25330 10362 25354 10364
rect 25410 10362 25434 10364
rect 25490 10362 25514 10364
rect 25570 10362 25576 10364
rect 25330 10310 25332 10362
rect 25512 10310 25514 10362
rect 25268 10308 25274 10310
rect 25330 10308 25354 10310
rect 25410 10308 25434 10310
rect 25490 10308 25514 10310
rect 25570 10308 25576 10310
rect 25268 10299 25576 10308
rect 21794 9820 22102 9829
rect 21794 9818 21800 9820
rect 21856 9818 21880 9820
rect 21936 9818 21960 9820
rect 22016 9818 22040 9820
rect 22096 9818 22102 9820
rect 21856 9766 21858 9818
rect 22038 9766 22040 9818
rect 21794 9764 21800 9766
rect 21856 9764 21880 9766
rect 21936 9764 21960 9766
rect 22016 9764 22040 9766
rect 22096 9764 22102 9766
rect 21794 9755 22102 9764
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 16684 7818 16712 9318
rect 18320 9276 18628 9285
rect 18320 9274 18326 9276
rect 18382 9274 18406 9276
rect 18462 9274 18486 9276
rect 18542 9274 18566 9276
rect 18622 9274 18628 9276
rect 18382 9222 18384 9274
rect 18564 9222 18566 9274
rect 18320 9220 18326 9222
rect 18382 9220 18406 9222
rect 18462 9220 18486 9222
rect 18542 9220 18566 9222
rect 18622 9220 18628 9222
rect 18320 9211 18628 9220
rect 18320 8188 18628 8197
rect 18320 8186 18326 8188
rect 18382 8186 18406 8188
rect 18462 8186 18486 8188
rect 18542 8186 18566 8188
rect 18622 8186 18628 8188
rect 18382 8134 18384 8186
rect 18564 8134 18566 8186
rect 18320 8132 18326 8134
rect 18382 8132 18406 8134
rect 18462 8132 18486 8134
rect 18542 8132 18566 8134
rect 18622 8132 18628 8134
rect 18320 8123 18628 8132
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 18320 7100 18628 7109
rect 18320 7098 18326 7100
rect 18382 7098 18406 7100
rect 18462 7098 18486 7100
rect 18542 7098 18566 7100
rect 18622 7098 18628 7100
rect 18382 7046 18384 7098
rect 18564 7046 18566 7098
rect 18320 7044 18326 7046
rect 18382 7044 18406 7046
rect 18462 7044 18486 7046
rect 18542 7044 18566 7046
rect 18622 7044 18628 7046
rect 18320 7035 18628 7044
rect 15212 6886 15332 6914
rect 15212 6798 15240 6886
rect 15200 6792 15252 6798
rect 18984 6769 19012 9318
rect 19628 9178 19656 9318
rect 25268 9276 25576 9285
rect 25268 9274 25274 9276
rect 25330 9274 25354 9276
rect 25410 9274 25434 9276
rect 25490 9274 25514 9276
rect 25570 9274 25576 9276
rect 25330 9222 25332 9274
rect 25512 9222 25514 9274
rect 25268 9220 25274 9222
rect 25330 9220 25354 9222
rect 25410 9220 25434 9222
rect 25490 9220 25514 9222
rect 25570 9220 25576 9222
rect 25268 9211 25576 9220
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 21794 8732 22102 8741
rect 21794 8730 21800 8732
rect 21856 8730 21880 8732
rect 21936 8730 21960 8732
rect 22016 8730 22040 8732
rect 22096 8730 22102 8732
rect 21856 8678 21858 8730
rect 22038 8678 22040 8730
rect 21794 8676 21800 8678
rect 21856 8676 21880 8678
rect 21936 8676 21960 8678
rect 22016 8676 22040 8678
rect 22096 8676 22102 8678
rect 21794 8667 22102 8676
rect 25268 8188 25576 8197
rect 25268 8186 25274 8188
rect 25330 8186 25354 8188
rect 25410 8186 25434 8188
rect 25490 8186 25514 8188
rect 25570 8186 25576 8188
rect 25330 8134 25332 8186
rect 25512 8134 25514 8186
rect 25268 8132 25274 8134
rect 25330 8132 25354 8134
rect 25410 8132 25434 8134
rect 25490 8132 25514 8134
rect 25570 8132 25576 8134
rect 25268 8123 25576 8132
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 21794 7644 22102 7653
rect 21794 7642 21800 7644
rect 21856 7642 21880 7644
rect 21936 7642 21960 7644
rect 22016 7642 22040 7644
rect 22096 7642 22102 7644
rect 21856 7590 21858 7642
rect 22038 7590 22040 7642
rect 21794 7588 21800 7590
rect 21856 7588 21880 7590
rect 21936 7588 21960 7590
rect 22016 7588 22040 7590
rect 22096 7588 22102 7590
rect 21794 7579 22102 7588
rect 15200 6734 15252 6740
rect 18970 6760 19026 6769
rect 14846 6556 15154 6565
rect 14846 6554 14852 6556
rect 14908 6554 14932 6556
rect 14988 6554 15012 6556
rect 15068 6554 15092 6556
rect 15148 6554 15154 6556
rect 14908 6502 14910 6554
rect 15090 6502 15092 6554
rect 14846 6500 14852 6502
rect 14908 6500 14932 6502
rect 14988 6500 15012 6502
rect 15068 6500 15092 6502
rect 15148 6500 15154 6502
rect 14846 6491 15154 6500
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14660 5234 14688 6394
rect 15212 6322 15240 6734
rect 18970 6695 19026 6704
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16592 6361 16620 6598
rect 21794 6556 22102 6565
rect 21794 6554 21800 6556
rect 21856 6554 21880 6556
rect 21936 6554 21960 6556
rect 22016 6554 22040 6556
rect 22096 6554 22102 6556
rect 21856 6502 21858 6554
rect 22038 6502 22040 6554
rect 21794 6500 21800 6502
rect 21856 6500 21880 6502
rect 21936 6500 21960 6502
rect 22016 6500 22040 6502
rect 22096 6500 22102 6502
rect 21794 6491 22102 6500
rect 16578 6352 16634 6361
rect 15200 6316 15252 6322
rect 16578 6287 16634 6296
rect 15200 6258 15252 6264
rect 15212 5710 15240 6258
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 10968 3120 11020 3126
rect 10968 3062 11020 3068
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 11992 2990 12020 3470
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14476 3194 14504 3402
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14752 3058 14780 5510
rect 14846 5468 15154 5477
rect 14846 5466 14852 5468
rect 14908 5466 14932 5468
rect 14988 5466 15012 5468
rect 15068 5466 15092 5468
rect 15148 5466 15154 5468
rect 14908 5414 14910 5466
rect 15090 5414 15092 5466
rect 14846 5412 14852 5414
rect 14908 5412 14932 5414
rect 14988 5412 15012 5414
rect 15068 5412 15092 5414
rect 15148 5412 15154 5414
rect 14846 5403 15154 5412
rect 16592 4826 16620 6287
rect 18320 6012 18628 6021
rect 18320 6010 18326 6012
rect 18382 6010 18406 6012
rect 18462 6010 18486 6012
rect 18542 6010 18566 6012
rect 18622 6010 18628 6012
rect 18382 5958 18384 6010
rect 18564 5958 18566 6010
rect 18320 5956 18326 5958
rect 18382 5956 18406 5958
rect 18462 5956 18486 5958
rect 18542 5956 18566 5958
rect 18622 5956 18628 5958
rect 18320 5947 18628 5956
rect 21794 5468 22102 5477
rect 21794 5466 21800 5468
rect 21856 5466 21880 5468
rect 21936 5466 21960 5468
rect 22016 5466 22040 5468
rect 22096 5466 22102 5468
rect 21856 5414 21858 5466
rect 22038 5414 22040 5466
rect 21794 5412 21800 5414
rect 21856 5412 21880 5414
rect 21936 5412 21960 5414
rect 22016 5412 22040 5414
rect 22096 5412 22102 5414
rect 21794 5403 22102 5412
rect 19892 5296 19944 5302
rect 19892 5238 19944 5244
rect 18320 4924 18628 4933
rect 18320 4922 18326 4924
rect 18382 4922 18406 4924
rect 18462 4922 18486 4924
rect 18542 4922 18566 4924
rect 18622 4922 18628 4924
rect 18382 4870 18384 4922
rect 18564 4870 18566 4922
rect 18320 4868 18326 4870
rect 18382 4868 18406 4870
rect 18462 4868 18486 4870
rect 18542 4868 18566 4870
rect 18622 4868 18628 4870
rect 18320 4859 18628 4868
rect 19904 4826 19932 5238
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 19892 4820 19944 4826
rect 19892 4762 19944 4768
rect 16592 4622 16620 4762
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16212 4548 16264 4554
rect 16212 4490 16264 4496
rect 14846 4380 15154 4389
rect 14846 4378 14852 4380
rect 14908 4378 14932 4380
rect 14988 4378 15012 4380
rect 15068 4378 15092 4380
rect 15148 4378 15154 4380
rect 14908 4326 14910 4378
rect 15090 4326 15092 4378
rect 14846 4324 14852 4326
rect 14908 4324 14932 4326
rect 14988 4324 15012 4326
rect 15068 4324 15092 4326
rect 15148 4324 15154 4326
rect 14846 4315 15154 4324
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 16132 3738 16160 4218
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16224 3534 16252 4490
rect 16396 4480 16448 4486
rect 16396 4422 16448 4428
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 14846 3292 15154 3301
rect 14846 3290 14852 3292
rect 14908 3290 14932 3292
rect 14988 3290 15012 3292
rect 15068 3290 15092 3292
rect 15148 3290 15154 3292
rect 14908 3238 14910 3290
rect 15090 3238 15092 3290
rect 14846 3236 14852 3238
rect 14908 3236 14932 3238
rect 14988 3236 15012 3238
rect 15068 3236 15092 3238
rect 15148 3236 15154 3238
rect 14846 3227 15154 3236
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 11372 2748 11680 2757
rect 11372 2746 11378 2748
rect 11434 2746 11458 2748
rect 11514 2746 11538 2748
rect 11594 2746 11618 2748
rect 11674 2746 11680 2748
rect 11434 2694 11436 2746
rect 11616 2694 11618 2746
rect 11372 2692 11378 2694
rect 11434 2692 11458 2694
rect 11514 2692 11538 2694
rect 11594 2692 11618 2694
rect 11674 2692 11680 2694
rect 11372 2683 11680 2692
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 16408 2378 16436 4422
rect 21794 4380 22102 4389
rect 21794 4378 21800 4380
rect 21856 4378 21880 4380
rect 21936 4378 21960 4380
rect 22016 4378 22040 4380
rect 22096 4378 22102 4380
rect 21856 4326 21858 4378
rect 22038 4326 22040 4378
rect 21794 4324 21800 4326
rect 21856 4324 21880 4326
rect 21936 4324 21960 4326
rect 22016 4324 22040 4326
rect 22096 4324 22102 4326
rect 21794 4315 22102 4324
rect 18320 3836 18628 3845
rect 18320 3834 18326 3836
rect 18382 3834 18406 3836
rect 18462 3834 18486 3836
rect 18542 3834 18566 3836
rect 18622 3834 18628 3836
rect 18382 3782 18384 3834
rect 18564 3782 18566 3834
rect 18320 3780 18326 3782
rect 18382 3780 18406 3782
rect 18462 3780 18486 3782
rect 18542 3780 18566 3782
rect 18622 3780 18628 3782
rect 18320 3771 18628 3780
rect 21794 3292 22102 3301
rect 21794 3290 21800 3292
rect 21856 3290 21880 3292
rect 21936 3290 21960 3292
rect 22016 3290 22040 3292
rect 22096 3290 22102 3292
rect 21856 3238 21858 3290
rect 22038 3238 22040 3290
rect 21794 3236 21800 3238
rect 21856 3236 21880 3238
rect 21936 3236 21960 3238
rect 22016 3236 22040 3238
rect 22096 3236 22102 3238
rect 21794 3227 22102 3236
rect 18320 2748 18628 2757
rect 18320 2746 18326 2748
rect 18382 2746 18406 2748
rect 18462 2746 18486 2748
rect 18542 2746 18566 2748
rect 18622 2746 18628 2748
rect 18382 2694 18384 2746
rect 18564 2694 18566 2746
rect 18320 2692 18326 2694
rect 18382 2692 18406 2694
rect 18462 2692 18486 2694
rect 18542 2692 18566 2694
rect 18622 2692 18628 2694
rect 18320 2683 18628 2692
rect 23308 2582 23336 7686
rect 25268 7100 25576 7109
rect 25268 7098 25274 7100
rect 25330 7098 25354 7100
rect 25410 7098 25434 7100
rect 25490 7098 25514 7100
rect 25570 7098 25576 7100
rect 25330 7046 25332 7098
rect 25512 7046 25514 7098
rect 25268 7044 25274 7046
rect 25330 7044 25354 7046
rect 25410 7044 25434 7046
rect 25490 7044 25514 7046
rect 25570 7044 25576 7046
rect 25268 7035 25576 7044
rect 25268 6012 25576 6021
rect 25268 6010 25274 6012
rect 25330 6010 25354 6012
rect 25410 6010 25434 6012
rect 25490 6010 25514 6012
rect 25570 6010 25576 6012
rect 25330 5958 25332 6010
rect 25512 5958 25514 6010
rect 25268 5956 25274 5958
rect 25330 5956 25354 5958
rect 25410 5956 25434 5958
rect 25490 5956 25514 5958
rect 25570 5956 25576 5958
rect 25268 5947 25576 5956
rect 25268 4924 25576 4933
rect 25268 4922 25274 4924
rect 25330 4922 25354 4924
rect 25410 4922 25434 4924
rect 25490 4922 25514 4924
rect 25570 4922 25576 4924
rect 25330 4870 25332 4922
rect 25512 4870 25514 4922
rect 25268 4868 25274 4870
rect 25330 4868 25354 4870
rect 25410 4868 25434 4870
rect 25490 4868 25514 4870
rect 25570 4868 25576 4870
rect 25268 4859 25576 4868
rect 25268 3836 25576 3845
rect 25268 3834 25274 3836
rect 25330 3834 25354 3836
rect 25410 3834 25434 3836
rect 25490 3834 25514 3836
rect 25570 3834 25576 3836
rect 25330 3782 25332 3834
rect 25512 3782 25514 3834
rect 25268 3780 25274 3782
rect 25330 3780 25354 3782
rect 25410 3780 25434 3782
rect 25490 3780 25514 3782
rect 25570 3780 25576 3782
rect 25268 3771 25576 3780
rect 25268 2748 25576 2757
rect 25268 2746 25274 2748
rect 25330 2746 25354 2748
rect 25410 2746 25434 2748
rect 25490 2746 25514 2748
rect 25570 2746 25576 2748
rect 25330 2694 25332 2746
rect 25512 2694 25514 2746
rect 25268 2692 25274 2694
rect 25330 2692 25354 2694
rect 25410 2692 25434 2694
rect 25490 2692 25514 2694
rect 25570 2692 25576 2694
rect 25268 2683 25576 2692
rect 23296 2576 23348 2582
rect 23296 2518 23348 2524
rect 2044 2372 2096 2378
rect 2044 2314 2096 2320
rect 16396 2372 16448 2378
rect 16396 2314 16448 2320
rect 23204 2372 23256 2378
rect 23204 2314 23256 2320
rect 7898 2204 8206 2213
rect 7898 2202 7904 2204
rect 7960 2202 7984 2204
rect 8040 2202 8064 2204
rect 8120 2202 8144 2204
rect 8200 2202 8206 2204
rect 7960 2150 7962 2202
rect 8142 2150 8144 2202
rect 7898 2148 7904 2150
rect 7960 2148 7984 2150
rect 8040 2148 8064 2150
rect 8120 2148 8144 2150
rect 8200 2148 8206 2150
rect 7898 2139 8206 2148
rect 14846 2204 15154 2213
rect 14846 2202 14852 2204
rect 14908 2202 14932 2204
rect 14988 2202 15012 2204
rect 15068 2202 15092 2204
rect 15148 2202 15154 2204
rect 14908 2150 14910 2202
rect 15090 2150 15092 2202
rect 14846 2148 14852 2150
rect 14908 2148 14932 2150
rect 14988 2148 15012 2150
rect 15068 2148 15092 2150
rect 15148 2148 15154 2150
rect 14846 2139 15154 2148
rect 21794 2204 22102 2213
rect 21794 2202 21800 2204
rect 21856 2202 21880 2204
rect 21936 2202 21960 2204
rect 22016 2202 22040 2204
rect 22096 2202 22102 2204
rect 21856 2150 21858 2202
rect 22038 2150 22040 2202
rect 21794 2148 21800 2150
rect 21856 2148 21880 2150
rect 21936 2148 21960 2150
rect 22016 2148 22040 2150
rect 22096 2148 22102 2150
rect 21794 2139 22102 2148
rect 23216 800 23244 2314
rect 18 0 74 800
rect 23202 0 23258 800
<< via2 >>
rect 4430 27770 4486 27772
rect 4510 27770 4566 27772
rect 4590 27770 4646 27772
rect 4670 27770 4726 27772
rect 4430 27718 4476 27770
rect 4476 27718 4486 27770
rect 4510 27718 4540 27770
rect 4540 27718 4552 27770
rect 4552 27718 4566 27770
rect 4590 27718 4604 27770
rect 4604 27718 4616 27770
rect 4616 27718 4646 27770
rect 4670 27718 4680 27770
rect 4680 27718 4726 27770
rect 4430 27716 4486 27718
rect 4510 27716 4566 27718
rect 4590 27716 4646 27718
rect 4670 27716 4726 27718
rect 11378 27770 11434 27772
rect 11458 27770 11514 27772
rect 11538 27770 11594 27772
rect 11618 27770 11674 27772
rect 11378 27718 11424 27770
rect 11424 27718 11434 27770
rect 11458 27718 11488 27770
rect 11488 27718 11500 27770
rect 11500 27718 11514 27770
rect 11538 27718 11552 27770
rect 11552 27718 11564 27770
rect 11564 27718 11594 27770
rect 11618 27718 11628 27770
rect 11628 27718 11674 27770
rect 11378 27716 11434 27718
rect 11458 27716 11514 27718
rect 11538 27716 11594 27718
rect 11618 27716 11674 27718
rect 18326 27770 18382 27772
rect 18406 27770 18462 27772
rect 18486 27770 18542 27772
rect 18566 27770 18622 27772
rect 18326 27718 18372 27770
rect 18372 27718 18382 27770
rect 18406 27718 18436 27770
rect 18436 27718 18448 27770
rect 18448 27718 18462 27770
rect 18486 27718 18500 27770
rect 18500 27718 18512 27770
rect 18512 27718 18542 27770
rect 18566 27718 18576 27770
rect 18576 27718 18622 27770
rect 18326 27716 18382 27718
rect 18406 27716 18462 27718
rect 18486 27716 18542 27718
rect 18566 27716 18622 27718
rect 25274 27770 25330 27772
rect 25354 27770 25410 27772
rect 25434 27770 25490 27772
rect 25514 27770 25570 27772
rect 25274 27718 25320 27770
rect 25320 27718 25330 27770
rect 25354 27718 25384 27770
rect 25384 27718 25396 27770
rect 25396 27718 25410 27770
rect 25434 27718 25448 27770
rect 25448 27718 25460 27770
rect 25460 27718 25490 27770
rect 25514 27718 25524 27770
rect 25524 27718 25570 27770
rect 25274 27716 25330 27718
rect 25354 27716 25410 27718
rect 25434 27716 25490 27718
rect 25514 27716 25570 27718
rect 7904 27226 7960 27228
rect 7984 27226 8040 27228
rect 8064 27226 8120 27228
rect 8144 27226 8200 27228
rect 7904 27174 7950 27226
rect 7950 27174 7960 27226
rect 7984 27174 8014 27226
rect 8014 27174 8026 27226
rect 8026 27174 8040 27226
rect 8064 27174 8078 27226
rect 8078 27174 8090 27226
rect 8090 27174 8120 27226
rect 8144 27174 8154 27226
rect 8154 27174 8200 27226
rect 7904 27172 7960 27174
rect 7984 27172 8040 27174
rect 8064 27172 8120 27174
rect 8144 27172 8200 27174
rect 14852 27226 14908 27228
rect 14932 27226 14988 27228
rect 15012 27226 15068 27228
rect 15092 27226 15148 27228
rect 14852 27174 14898 27226
rect 14898 27174 14908 27226
rect 14932 27174 14962 27226
rect 14962 27174 14974 27226
rect 14974 27174 14988 27226
rect 15012 27174 15026 27226
rect 15026 27174 15038 27226
rect 15038 27174 15068 27226
rect 15092 27174 15102 27226
rect 15102 27174 15148 27226
rect 14852 27172 14908 27174
rect 14932 27172 14988 27174
rect 15012 27172 15068 27174
rect 15092 27172 15148 27174
rect 4430 26682 4486 26684
rect 4510 26682 4566 26684
rect 4590 26682 4646 26684
rect 4670 26682 4726 26684
rect 4430 26630 4476 26682
rect 4476 26630 4486 26682
rect 4510 26630 4540 26682
rect 4540 26630 4552 26682
rect 4552 26630 4566 26682
rect 4590 26630 4604 26682
rect 4604 26630 4616 26682
rect 4616 26630 4646 26682
rect 4670 26630 4680 26682
rect 4680 26630 4726 26682
rect 4430 26628 4486 26630
rect 4510 26628 4566 26630
rect 4590 26628 4646 26630
rect 4670 26628 4726 26630
rect 11378 26682 11434 26684
rect 11458 26682 11514 26684
rect 11538 26682 11594 26684
rect 11618 26682 11674 26684
rect 11378 26630 11424 26682
rect 11424 26630 11434 26682
rect 11458 26630 11488 26682
rect 11488 26630 11500 26682
rect 11500 26630 11514 26682
rect 11538 26630 11552 26682
rect 11552 26630 11564 26682
rect 11564 26630 11594 26682
rect 11618 26630 11628 26682
rect 11628 26630 11674 26682
rect 11378 26628 11434 26630
rect 11458 26628 11514 26630
rect 11538 26628 11594 26630
rect 11618 26628 11674 26630
rect 7904 26138 7960 26140
rect 7984 26138 8040 26140
rect 8064 26138 8120 26140
rect 8144 26138 8200 26140
rect 7904 26086 7950 26138
rect 7950 26086 7960 26138
rect 7984 26086 8014 26138
rect 8014 26086 8026 26138
rect 8026 26086 8040 26138
rect 8064 26086 8078 26138
rect 8078 26086 8090 26138
rect 8090 26086 8120 26138
rect 8144 26086 8154 26138
rect 8154 26086 8200 26138
rect 7904 26084 7960 26086
rect 7984 26084 8040 26086
rect 8064 26084 8120 26086
rect 8144 26084 8200 26086
rect 14852 26138 14908 26140
rect 14932 26138 14988 26140
rect 15012 26138 15068 26140
rect 15092 26138 15148 26140
rect 14852 26086 14898 26138
rect 14898 26086 14908 26138
rect 14932 26086 14962 26138
rect 14962 26086 14974 26138
rect 14974 26086 14988 26138
rect 15012 26086 15026 26138
rect 15026 26086 15038 26138
rect 15038 26086 15068 26138
rect 15092 26086 15102 26138
rect 15102 26086 15148 26138
rect 14852 26084 14908 26086
rect 14932 26084 14988 26086
rect 15012 26084 15068 26086
rect 15092 26084 15148 26086
rect 4430 25594 4486 25596
rect 4510 25594 4566 25596
rect 4590 25594 4646 25596
rect 4670 25594 4726 25596
rect 4430 25542 4476 25594
rect 4476 25542 4486 25594
rect 4510 25542 4540 25594
rect 4540 25542 4552 25594
rect 4552 25542 4566 25594
rect 4590 25542 4604 25594
rect 4604 25542 4616 25594
rect 4616 25542 4646 25594
rect 4670 25542 4680 25594
rect 4680 25542 4726 25594
rect 4430 25540 4486 25542
rect 4510 25540 4566 25542
rect 4590 25540 4646 25542
rect 4670 25540 4726 25542
rect 11378 25594 11434 25596
rect 11458 25594 11514 25596
rect 11538 25594 11594 25596
rect 11618 25594 11674 25596
rect 11378 25542 11424 25594
rect 11424 25542 11434 25594
rect 11458 25542 11488 25594
rect 11488 25542 11500 25594
rect 11500 25542 11514 25594
rect 11538 25542 11552 25594
rect 11552 25542 11564 25594
rect 11564 25542 11594 25594
rect 11618 25542 11628 25594
rect 11628 25542 11674 25594
rect 11378 25540 11434 25542
rect 11458 25540 11514 25542
rect 11538 25540 11594 25542
rect 11618 25540 11674 25542
rect 7904 25050 7960 25052
rect 7984 25050 8040 25052
rect 8064 25050 8120 25052
rect 8144 25050 8200 25052
rect 7904 24998 7950 25050
rect 7950 24998 7960 25050
rect 7984 24998 8014 25050
rect 8014 24998 8026 25050
rect 8026 24998 8040 25050
rect 8064 24998 8078 25050
rect 8078 24998 8090 25050
rect 8090 24998 8120 25050
rect 8144 24998 8154 25050
rect 8154 24998 8200 25050
rect 7904 24996 7960 24998
rect 7984 24996 8040 24998
rect 8064 24996 8120 24998
rect 8144 24996 8200 24998
rect 14852 25050 14908 25052
rect 14932 25050 14988 25052
rect 15012 25050 15068 25052
rect 15092 25050 15148 25052
rect 14852 24998 14898 25050
rect 14898 24998 14908 25050
rect 14932 24998 14962 25050
rect 14962 24998 14974 25050
rect 14974 24998 14988 25050
rect 15012 24998 15026 25050
rect 15026 24998 15038 25050
rect 15038 24998 15068 25050
rect 15092 24998 15102 25050
rect 15102 24998 15148 25050
rect 14852 24996 14908 24998
rect 14932 24996 14988 24998
rect 15012 24996 15068 24998
rect 15092 24996 15148 24998
rect 1490 24556 1492 24576
rect 1492 24556 1544 24576
rect 1544 24556 1546 24576
rect 1490 24520 1546 24556
rect 4430 24506 4486 24508
rect 4510 24506 4566 24508
rect 4590 24506 4646 24508
rect 4670 24506 4726 24508
rect 4430 24454 4476 24506
rect 4476 24454 4486 24506
rect 4510 24454 4540 24506
rect 4540 24454 4552 24506
rect 4552 24454 4566 24506
rect 4590 24454 4604 24506
rect 4604 24454 4616 24506
rect 4616 24454 4646 24506
rect 4670 24454 4680 24506
rect 4680 24454 4726 24506
rect 4430 24452 4486 24454
rect 4510 24452 4566 24454
rect 4590 24452 4646 24454
rect 4670 24452 4726 24454
rect 4430 23418 4486 23420
rect 4510 23418 4566 23420
rect 4590 23418 4646 23420
rect 4670 23418 4726 23420
rect 4430 23366 4476 23418
rect 4476 23366 4486 23418
rect 4510 23366 4540 23418
rect 4540 23366 4552 23418
rect 4552 23366 4566 23418
rect 4590 23366 4604 23418
rect 4604 23366 4616 23418
rect 4616 23366 4646 23418
rect 4670 23366 4680 23418
rect 4680 23366 4726 23418
rect 4430 23364 4486 23366
rect 4510 23364 4566 23366
rect 4590 23364 4646 23366
rect 4670 23364 4726 23366
rect 4430 22330 4486 22332
rect 4510 22330 4566 22332
rect 4590 22330 4646 22332
rect 4670 22330 4726 22332
rect 4430 22278 4476 22330
rect 4476 22278 4486 22330
rect 4510 22278 4540 22330
rect 4540 22278 4552 22330
rect 4552 22278 4566 22330
rect 4590 22278 4604 22330
rect 4604 22278 4616 22330
rect 4616 22278 4646 22330
rect 4670 22278 4680 22330
rect 4680 22278 4726 22330
rect 4430 22276 4486 22278
rect 4510 22276 4566 22278
rect 4590 22276 4646 22278
rect 4670 22276 4726 22278
rect 4430 21242 4486 21244
rect 4510 21242 4566 21244
rect 4590 21242 4646 21244
rect 4670 21242 4726 21244
rect 4430 21190 4476 21242
rect 4476 21190 4486 21242
rect 4510 21190 4540 21242
rect 4540 21190 4552 21242
rect 4552 21190 4566 21242
rect 4590 21190 4604 21242
rect 4604 21190 4616 21242
rect 4616 21190 4646 21242
rect 4670 21190 4680 21242
rect 4680 21190 4726 21242
rect 4430 21188 4486 21190
rect 4510 21188 4566 21190
rect 4590 21188 4646 21190
rect 4670 21188 4726 21190
rect 4430 20154 4486 20156
rect 4510 20154 4566 20156
rect 4590 20154 4646 20156
rect 4670 20154 4726 20156
rect 4430 20102 4476 20154
rect 4476 20102 4486 20154
rect 4510 20102 4540 20154
rect 4540 20102 4552 20154
rect 4552 20102 4566 20154
rect 4590 20102 4604 20154
rect 4604 20102 4616 20154
rect 4616 20102 4646 20154
rect 4670 20102 4680 20154
rect 4680 20102 4726 20154
rect 4430 20100 4486 20102
rect 4510 20100 4566 20102
rect 4590 20100 4646 20102
rect 4670 20100 4726 20102
rect 4430 19066 4486 19068
rect 4510 19066 4566 19068
rect 4590 19066 4646 19068
rect 4670 19066 4726 19068
rect 4430 19014 4476 19066
rect 4476 19014 4486 19066
rect 4510 19014 4540 19066
rect 4540 19014 4552 19066
rect 4552 19014 4566 19066
rect 4590 19014 4604 19066
rect 4604 19014 4616 19066
rect 4616 19014 4646 19066
rect 4670 19014 4680 19066
rect 4680 19014 4726 19066
rect 4430 19012 4486 19014
rect 4510 19012 4566 19014
rect 4590 19012 4646 19014
rect 4670 19012 4726 19014
rect 4430 17978 4486 17980
rect 4510 17978 4566 17980
rect 4590 17978 4646 17980
rect 4670 17978 4726 17980
rect 4430 17926 4476 17978
rect 4476 17926 4486 17978
rect 4510 17926 4540 17978
rect 4540 17926 4552 17978
rect 4552 17926 4566 17978
rect 4590 17926 4604 17978
rect 4604 17926 4616 17978
rect 4616 17926 4646 17978
rect 4670 17926 4680 17978
rect 4680 17926 4726 17978
rect 4430 17924 4486 17926
rect 4510 17924 4566 17926
rect 4590 17924 4646 17926
rect 4670 17924 4726 17926
rect 4430 16890 4486 16892
rect 4510 16890 4566 16892
rect 4590 16890 4646 16892
rect 4670 16890 4726 16892
rect 4430 16838 4476 16890
rect 4476 16838 4486 16890
rect 4510 16838 4540 16890
rect 4540 16838 4552 16890
rect 4552 16838 4566 16890
rect 4590 16838 4604 16890
rect 4604 16838 4616 16890
rect 4616 16838 4646 16890
rect 4670 16838 4680 16890
rect 4680 16838 4726 16890
rect 4430 16836 4486 16838
rect 4510 16836 4566 16838
rect 4590 16836 4646 16838
rect 4670 16836 4726 16838
rect 4430 15802 4486 15804
rect 4510 15802 4566 15804
rect 4590 15802 4646 15804
rect 4670 15802 4726 15804
rect 4430 15750 4476 15802
rect 4476 15750 4486 15802
rect 4510 15750 4540 15802
rect 4540 15750 4552 15802
rect 4552 15750 4566 15802
rect 4590 15750 4604 15802
rect 4604 15750 4616 15802
rect 4616 15750 4646 15802
rect 4670 15750 4680 15802
rect 4680 15750 4726 15802
rect 4430 15748 4486 15750
rect 4510 15748 4566 15750
rect 4590 15748 4646 15750
rect 4670 15748 4726 15750
rect 11378 24506 11434 24508
rect 11458 24506 11514 24508
rect 11538 24506 11594 24508
rect 11618 24506 11674 24508
rect 11378 24454 11424 24506
rect 11424 24454 11434 24506
rect 11458 24454 11488 24506
rect 11488 24454 11500 24506
rect 11500 24454 11514 24506
rect 11538 24454 11552 24506
rect 11552 24454 11564 24506
rect 11564 24454 11594 24506
rect 11618 24454 11628 24506
rect 11628 24454 11674 24506
rect 11378 24452 11434 24454
rect 11458 24452 11514 24454
rect 11538 24452 11594 24454
rect 11618 24452 11674 24454
rect 7904 23962 7960 23964
rect 7984 23962 8040 23964
rect 8064 23962 8120 23964
rect 8144 23962 8200 23964
rect 7904 23910 7950 23962
rect 7950 23910 7960 23962
rect 7984 23910 8014 23962
rect 8014 23910 8026 23962
rect 8026 23910 8040 23962
rect 8064 23910 8078 23962
rect 8078 23910 8090 23962
rect 8090 23910 8120 23962
rect 8144 23910 8154 23962
rect 8154 23910 8200 23962
rect 7904 23908 7960 23910
rect 7984 23908 8040 23910
rect 8064 23908 8120 23910
rect 8144 23908 8200 23910
rect 14852 23962 14908 23964
rect 14932 23962 14988 23964
rect 15012 23962 15068 23964
rect 15092 23962 15148 23964
rect 14852 23910 14898 23962
rect 14898 23910 14908 23962
rect 14932 23910 14962 23962
rect 14962 23910 14974 23962
rect 14974 23910 14988 23962
rect 15012 23910 15026 23962
rect 15026 23910 15038 23962
rect 15038 23910 15068 23962
rect 15092 23910 15102 23962
rect 15102 23910 15148 23962
rect 14852 23908 14908 23910
rect 14932 23908 14988 23910
rect 15012 23908 15068 23910
rect 15092 23908 15148 23910
rect 11378 23418 11434 23420
rect 11458 23418 11514 23420
rect 11538 23418 11594 23420
rect 11618 23418 11674 23420
rect 11378 23366 11424 23418
rect 11424 23366 11434 23418
rect 11458 23366 11488 23418
rect 11488 23366 11500 23418
rect 11500 23366 11514 23418
rect 11538 23366 11552 23418
rect 11552 23366 11564 23418
rect 11564 23366 11594 23418
rect 11618 23366 11628 23418
rect 11628 23366 11674 23418
rect 11378 23364 11434 23366
rect 11458 23364 11514 23366
rect 11538 23364 11594 23366
rect 11618 23364 11674 23366
rect 7904 22874 7960 22876
rect 7984 22874 8040 22876
rect 8064 22874 8120 22876
rect 8144 22874 8200 22876
rect 7904 22822 7950 22874
rect 7950 22822 7960 22874
rect 7984 22822 8014 22874
rect 8014 22822 8026 22874
rect 8026 22822 8040 22874
rect 8064 22822 8078 22874
rect 8078 22822 8090 22874
rect 8090 22822 8120 22874
rect 8144 22822 8154 22874
rect 8154 22822 8200 22874
rect 7904 22820 7960 22822
rect 7984 22820 8040 22822
rect 8064 22820 8120 22822
rect 8144 22820 8200 22822
rect 14852 22874 14908 22876
rect 14932 22874 14988 22876
rect 15012 22874 15068 22876
rect 15092 22874 15148 22876
rect 14852 22822 14898 22874
rect 14898 22822 14908 22874
rect 14932 22822 14962 22874
rect 14962 22822 14974 22874
rect 14974 22822 14988 22874
rect 15012 22822 15026 22874
rect 15026 22822 15038 22874
rect 15038 22822 15068 22874
rect 15092 22822 15102 22874
rect 15102 22822 15148 22874
rect 14852 22820 14908 22822
rect 14932 22820 14988 22822
rect 15012 22820 15068 22822
rect 15092 22820 15148 22822
rect 11378 22330 11434 22332
rect 11458 22330 11514 22332
rect 11538 22330 11594 22332
rect 11618 22330 11674 22332
rect 11378 22278 11424 22330
rect 11424 22278 11434 22330
rect 11458 22278 11488 22330
rect 11488 22278 11500 22330
rect 11500 22278 11514 22330
rect 11538 22278 11552 22330
rect 11552 22278 11564 22330
rect 11564 22278 11594 22330
rect 11618 22278 11628 22330
rect 11628 22278 11674 22330
rect 11378 22276 11434 22278
rect 11458 22276 11514 22278
rect 11538 22276 11594 22278
rect 11618 22276 11674 22278
rect 7904 21786 7960 21788
rect 7984 21786 8040 21788
rect 8064 21786 8120 21788
rect 8144 21786 8200 21788
rect 7904 21734 7950 21786
rect 7950 21734 7960 21786
rect 7984 21734 8014 21786
rect 8014 21734 8026 21786
rect 8026 21734 8040 21786
rect 8064 21734 8078 21786
rect 8078 21734 8090 21786
rect 8090 21734 8120 21786
rect 8144 21734 8154 21786
rect 8154 21734 8200 21786
rect 7904 21732 7960 21734
rect 7984 21732 8040 21734
rect 8064 21732 8120 21734
rect 8144 21732 8200 21734
rect 14852 21786 14908 21788
rect 14932 21786 14988 21788
rect 15012 21786 15068 21788
rect 15092 21786 15148 21788
rect 14852 21734 14898 21786
rect 14898 21734 14908 21786
rect 14932 21734 14962 21786
rect 14962 21734 14974 21786
rect 14974 21734 14988 21786
rect 15012 21734 15026 21786
rect 15026 21734 15038 21786
rect 15038 21734 15068 21786
rect 15092 21734 15102 21786
rect 15102 21734 15148 21786
rect 14852 21732 14908 21734
rect 14932 21732 14988 21734
rect 15012 21732 15068 21734
rect 15092 21732 15148 21734
rect 11378 21242 11434 21244
rect 11458 21242 11514 21244
rect 11538 21242 11594 21244
rect 11618 21242 11674 21244
rect 11378 21190 11424 21242
rect 11424 21190 11434 21242
rect 11458 21190 11488 21242
rect 11488 21190 11500 21242
rect 11500 21190 11514 21242
rect 11538 21190 11552 21242
rect 11552 21190 11564 21242
rect 11564 21190 11594 21242
rect 11618 21190 11628 21242
rect 11628 21190 11674 21242
rect 11378 21188 11434 21190
rect 11458 21188 11514 21190
rect 11538 21188 11594 21190
rect 11618 21188 11674 21190
rect 7904 20698 7960 20700
rect 7984 20698 8040 20700
rect 8064 20698 8120 20700
rect 8144 20698 8200 20700
rect 7904 20646 7950 20698
rect 7950 20646 7960 20698
rect 7984 20646 8014 20698
rect 8014 20646 8026 20698
rect 8026 20646 8040 20698
rect 8064 20646 8078 20698
rect 8078 20646 8090 20698
rect 8090 20646 8120 20698
rect 8144 20646 8154 20698
rect 8154 20646 8200 20698
rect 7904 20644 7960 20646
rect 7984 20644 8040 20646
rect 8064 20644 8120 20646
rect 8144 20644 8200 20646
rect 14852 20698 14908 20700
rect 14932 20698 14988 20700
rect 15012 20698 15068 20700
rect 15092 20698 15148 20700
rect 14852 20646 14898 20698
rect 14898 20646 14908 20698
rect 14932 20646 14962 20698
rect 14962 20646 14974 20698
rect 14974 20646 14988 20698
rect 15012 20646 15026 20698
rect 15026 20646 15038 20698
rect 15038 20646 15068 20698
rect 15092 20646 15102 20698
rect 15102 20646 15148 20698
rect 14852 20644 14908 20646
rect 14932 20644 14988 20646
rect 15012 20644 15068 20646
rect 15092 20644 15148 20646
rect 11378 20154 11434 20156
rect 11458 20154 11514 20156
rect 11538 20154 11594 20156
rect 11618 20154 11674 20156
rect 11378 20102 11424 20154
rect 11424 20102 11434 20154
rect 11458 20102 11488 20154
rect 11488 20102 11500 20154
rect 11500 20102 11514 20154
rect 11538 20102 11552 20154
rect 11552 20102 11564 20154
rect 11564 20102 11594 20154
rect 11618 20102 11628 20154
rect 11628 20102 11674 20154
rect 11378 20100 11434 20102
rect 11458 20100 11514 20102
rect 11538 20100 11594 20102
rect 11618 20100 11674 20102
rect 7904 19610 7960 19612
rect 7984 19610 8040 19612
rect 8064 19610 8120 19612
rect 8144 19610 8200 19612
rect 7904 19558 7950 19610
rect 7950 19558 7960 19610
rect 7984 19558 8014 19610
rect 8014 19558 8026 19610
rect 8026 19558 8040 19610
rect 8064 19558 8078 19610
rect 8078 19558 8090 19610
rect 8090 19558 8120 19610
rect 8144 19558 8154 19610
rect 8154 19558 8200 19610
rect 7904 19556 7960 19558
rect 7984 19556 8040 19558
rect 8064 19556 8120 19558
rect 8144 19556 8200 19558
rect 14852 19610 14908 19612
rect 14932 19610 14988 19612
rect 15012 19610 15068 19612
rect 15092 19610 15148 19612
rect 14852 19558 14898 19610
rect 14898 19558 14908 19610
rect 14932 19558 14962 19610
rect 14962 19558 14974 19610
rect 14974 19558 14988 19610
rect 15012 19558 15026 19610
rect 15026 19558 15038 19610
rect 15038 19558 15068 19610
rect 15092 19558 15102 19610
rect 15102 19558 15148 19610
rect 14852 19556 14908 19558
rect 14932 19556 14988 19558
rect 15012 19556 15068 19558
rect 15092 19556 15148 19558
rect 11378 19066 11434 19068
rect 11458 19066 11514 19068
rect 11538 19066 11594 19068
rect 11618 19066 11674 19068
rect 11378 19014 11424 19066
rect 11424 19014 11434 19066
rect 11458 19014 11488 19066
rect 11488 19014 11500 19066
rect 11500 19014 11514 19066
rect 11538 19014 11552 19066
rect 11552 19014 11564 19066
rect 11564 19014 11594 19066
rect 11618 19014 11628 19066
rect 11628 19014 11674 19066
rect 11378 19012 11434 19014
rect 11458 19012 11514 19014
rect 11538 19012 11594 19014
rect 11618 19012 11674 19014
rect 7904 18522 7960 18524
rect 7984 18522 8040 18524
rect 8064 18522 8120 18524
rect 8144 18522 8200 18524
rect 7904 18470 7950 18522
rect 7950 18470 7960 18522
rect 7984 18470 8014 18522
rect 8014 18470 8026 18522
rect 8026 18470 8040 18522
rect 8064 18470 8078 18522
rect 8078 18470 8090 18522
rect 8090 18470 8120 18522
rect 8144 18470 8154 18522
rect 8154 18470 8200 18522
rect 7904 18468 7960 18470
rect 7984 18468 8040 18470
rect 8064 18468 8120 18470
rect 8144 18468 8200 18470
rect 14852 18522 14908 18524
rect 14932 18522 14988 18524
rect 15012 18522 15068 18524
rect 15092 18522 15148 18524
rect 14852 18470 14898 18522
rect 14898 18470 14908 18522
rect 14932 18470 14962 18522
rect 14962 18470 14974 18522
rect 14974 18470 14988 18522
rect 15012 18470 15026 18522
rect 15026 18470 15038 18522
rect 15038 18470 15068 18522
rect 15092 18470 15102 18522
rect 15102 18470 15148 18522
rect 14852 18468 14908 18470
rect 14932 18468 14988 18470
rect 15012 18468 15068 18470
rect 15092 18468 15148 18470
rect 11378 17978 11434 17980
rect 11458 17978 11514 17980
rect 11538 17978 11594 17980
rect 11618 17978 11674 17980
rect 11378 17926 11424 17978
rect 11424 17926 11434 17978
rect 11458 17926 11488 17978
rect 11488 17926 11500 17978
rect 11500 17926 11514 17978
rect 11538 17926 11552 17978
rect 11552 17926 11564 17978
rect 11564 17926 11594 17978
rect 11618 17926 11628 17978
rect 11628 17926 11674 17978
rect 11378 17924 11434 17926
rect 11458 17924 11514 17926
rect 11538 17924 11594 17926
rect 11618 17924 11674 17926
rect 7904 17434 7960 17436
rect 7984 17434 8040 17436
rect 8064 17434 8120 17436
rect 8144 17434 8200 17436
rect 7904 17382 7950 17434
rect 7950 17382 7960 17434
rect 7984 17382 8014 17434
rect 8014 17382 8026 17434
rect 8026 17382 8040 17434
rect 8064 17382 8078 17434
rect 8078 17382 8090 17434
rect 8090 17382 8120 17434
rect 8144 17382 8154 17434
rect 8154 17382 8200 17434
rect 7904 17380 7960 17382
rect 7984 17380 8040 17382
rect 8064 17380 8120 17382
rect 8144 17380 8200 17382
rect 14852 17434 14908 17436
rect 14932 17434 14988 17436
rect 15012 17434 15068 17436
rect 15092 17434 15148 17436
rect 14852 17382 14898 17434
rect 14898 17382 14908 17434
rect 14932 17382 14962 17434
rect 14962 17382 14974 17434
rect 14974 17382 14988 17434
rect 15012 17382 15026 17434
rect 15026 17382 15038 17434
rect 15038 17382 15068 17434
rect 15092 17382 15102 17434
rect 15102 17382 15148 17434
rect 14852 17380 14908 17382
rect 14932 17380 14988 17382
rect 15012 17380 15068 17382
rect 15092 17380 15148 17382
rect 4430 14714 4486 14716
rect 4510 14714 4566 14716
rect 4590 14714 4646 14716
rect 4670 14714 4726 14716
rect 4430 14662 4476 14714
rect 4476 14662 4486 14714
rect 4510 14662 4540 14714
rect 4540 14662 4552 14714
rect 4552 14662 4566 14714
rect 4590 14662 4604 14714
rect 4604 14662 4616 14714
rect 4616 14662 4646 14714
rect 4670 14662 4680 14714
rect 4680 14662 4726 14714
rect 4430 14660 4486 14662
rect 4510 14660 4566 14662
rect 4590 14660 4646 14662
rect 4670 14660 4726 14662
rect 4430 13626 4486 13628
rect 4510 13626 4566 13628
rect 4590 13626 4646 13628
rect 4670 13626 4726 13628
rect 4430 13574 4476 13626
rect 4476 13574 4486 13626
rect 4510 13574 4540 13626
rect 4540 13574 4552 13626
rect 4552 13574 4566 13626
rect 4590 13574 4604 13626
rect 4604 13574 4616 13626
rect 4616 13574 4646 13626
rect 4670 13574 4680 13626
rect 4680 13574 4726 13626
rect 4430 13572 4486 13574
rect 4510 13572 4566 13574
rect 4590 13572 4646 13574
rect 4670 13572 4726 13574
rect 4250 13252 4306 13288
rect 4250 13232 4252 13252
rect 4252 13232 4304 13252
rect 4304 13232 4306 13252
rect 4430 12538 4486 12540
rect 4510 12538 4566 12540
rect 4590 12538 4646 12540
rect 4670 12538 4726 12540
rect 4430 12486 4476 12538
rect 4476 12486 4486 12538
rect 4510 12486 4540 12538
rect 4540 12486 4552 12538
rect 4552 12486 4566 12538
rect 4590 12486 4604 12538
rect 4604 12486 4616 12538
rect 4616 12486 4646 12538
rect 4670 12486 4680 12538
rect 4680 12486 4726 12538
rect 4430 12484 4486 12486
rect 4510 12484 4566 12486
rect 4590 12484 4646 12486
rect 4670 12484 4726 12486
rect 4430 11450 4486 11452
rect 4510 11450 4566 11452
rect 4590 11450 4646 11452
rect 4670 11450 4726 11452
rect 4430 11398 4476 11450
rect 4476 11398 4486 11450
rect 4510 11398 4540 11450
rect 4540 11398 4552 11450
rect 4552 11398 4566 11450
rect 4590 11398 4604 11450
rect 4604 11398 4616 11450
rect 4616 11398 4646 11450
rect 4670 11398 4680 11450
rect 4680 11398 4726 11450
rect 4430 11396 4486 11398
rect 4510 11396 4566 11398
rect 4590 11396 4646 11398
rect 4670 11396 4726 11398
rect 4430 10362 4486 10364
rect 4510 10362 4566 10364
rect 4590 10362 4646 10364
rect 4670 10362 4726 10364
rect 4430 10310 4476 10362
rect 4476 10310 4486 10362
rect 4510 10310 4540 10362
rect 4540 10310 4552 10362
rect 4552 10310 4566 10362
rect 4590 10310 4604 10362
rect 4604 10310 4616 10362
rect 4616 10310 4646 10362
rect 4670 10310 4680 10362
rect 4680 10310 4726 10362
rect 4430 10308 4486 10310
rect 4510 10308 4566 10310
rect 4590 10308 4646 10310
rect 4670 10308 4726 10310
rect 4430 9274 4486 9276
rect 4510 9274 4566 9276
rect 4590 9274 4646 9276
rect 4670 9274 4726 9276
rect 4430 9222 4476 9274
rect 4476 9222 4486 9274
rect 4510 9222 4540 9274
rect 4540 9222 4552 9274
rect 4552 9222 4566 9274
rect 4590 9222 4604 9274
rect 4604 9222 4616 9274
rect 4616 9222 4646 9274
rect 4670 9222 4680 9274
rect 4680 9222 4726 9274
rect 4430 9220 4486 9222
rect 4510 9220 4566 9222
rect 4590 9220 4646 9222
rect 4670 9220 4726 9222
rect 7904 16346 7960 16348
rect 7984 16346 8040 16348
rect 8064 16346 8120 16348
rect 8144 16346 8200 16348
rect 7904 16294 7950 16346
rect 7950 16294 7960 16346
rect 7984 16294 8014 16346
rect 8014 16294 8026 16346
rect 8026 16294 8040 16346
rect 8064 16294 8078 16346
rect 8078 16294 8090 16346
rect 8090 16294 8120 16346
rect 8144 16294 8154 16346
rect 8154 16294 8200 16346
rect 7904 16292 7960 16294
rect 7984 16292 8040 16294
rect 8064 16292 8120 16294
rect 8144 16292 8200 16294
rect 11378 16890 11434 16892
rect 11458 16890 11514 16892
rect 11538 16890 11594 16892
rect 11618 16890 11674 16892
rect 11378 16838 11424 16890
rect 11424 16838 11434 16890
rect 11458 16838 11488 16890
rect 11488 16838 11500 16890
rect 11500 16838 11514 16890
rect 11538 16838 11552 16890
rect 11552 16838 11564 16890
rect 11564 16838 11594 16890
rect 11618 16838 11628 16890
rect 11628 16838 11674 16890
rect 11378 16836 11434 16838
rect 11458 16836 11514 16838
rect 11538 16836 11594 16838
rect 11618 16836 11674 16838
rect 7904 15258 7960 15260
rect 7984 15258 8040 15260
rect 8064 15258 8120 15260
rect 8144 15258 8200 15260
rect 7904 15206 7950 15258
rect 7950 15206 7960 15258
rect 7984 15206 8014 15258
rect 8014 15206 8026 15258
rect 8026 15206 8040 15258
rect 8064 15206 8078 15258
rect 8078 15206 8090 15258
rect 8090 15206 8120 15258
rect 8144 15206 8154 15258
rect 8154 15206 8200 15258
rect 7904 15204 7960 15206
rect 7984 15204 8040 15206
rect 8064 15204 8120 15206
rect 8144 15204 8200 15206
rect 7904 14170 7960 14172
rect 7984 14170 8040 14172
rect 8064 14170 8120 14172
rect 8144 14170 8200 14172
rect 7904 14118 7950 14170
rect 7950 14118 7960 14170
rect 7984 14118 8014 14170
rect 8014 14118 8026 14170
rect 8026 14118 8040 14170
rect 8064 14118 8078 14170
rect 8078 14118 8090 14170
rect 8090 14118 8120 14170
rect 8144 14118 8154 14170
rect 8154 14118 8200 14170
rect 7904 14116 7960 14118
rect 7984 14116 8040 14118
rect 8064 14116 8120 14118
rect 8144 14116 8200 14118
rect 4430 8186 4486 8188
rect 4510 8186 4566 8188
rect 4590 8186 4646 8188
rect 4670 8186 4726 8188
rect 4430 8134 4476 8186
rect 4476 8134 4486 8186
rect 4510 8134 4540 8186
rect 4540 8134 4552 8186
rect 4552 8134 4566 8186
rect 4590 8134 4604 8186
rect 4604 8134 4616 8186
rect 4616 8134 4646 8186
rect 4670 8134 4680 8186
rect 4680 8134 4726 8186
rect 4430 8132 4486 8134
rect 4510 8132 4566 8134
rect 4590 8132 4646 8134
rect 4670 8132 4726 8134
rect 4430 7098 4486 7100
rect 4510 7098 4566 7100
rect 4590 7098 4646 7100
rect 4670 7098 4726 7100
rect 4430 7046 4476 7098
rect 4476 7046 4486 7098
rect 4510 7046 4540 7098
rect 4540 7046 4552 7098
rect 4552 7046 4566 7098
rect 4590 7046 4604 7098
rect 4604 7046 4616 7098
rect 4616 7046 4646 7098
rect 4670 7046 4680 7098
rect 4680 7046 4726 7098
rect 4430 7044 4486 7046
rect 4510 7044 4566 7046
rect 4590 7044 4646 7046
rect 4670 7044 4726 7046
rect 4430 6010 4486 6012
rect 4510 6010 4566 6012
rect 4590 6010 4646 6012
rect 4670 6010 4726 6012
rect 4430 5958 4476 6010
rect 4476 5958 4486 6010
rect 4510 5958 4540 6010
rect 4540 5958 4552 6010
rect 4552 5958 4566 6010
rect 4590 5958 4604 6010
rect 4604 5958 4616 6010
rect 4616 5958 4646 6010
rect 4670 5958 4680 6010
rect 4680 5958 4726 6010
rect 4430 5956 4486 5958
rect 4510 5956 4566 5958
rect 4590 5956 4646 5958
rect 4670 5956 4726 5958
rect 5906 6840 5962 6896
rect 5354 6332 5356 6352
rect 5356 6332 5408 6352
rect 5408 6332 5410 6352
rect 5354 6296 5410 6332
rect 4430 4922 4486 4924
rect 4510 4922 4566 4924
rect 4590 4922 4646 4924
rect 4670 4922 4726 4924
rect 4430 4870 4476 4922
rect 4476 4870 4486 4922
rect 4510 4870 4540 4922
rect 4540 4870 4552 4922
rect 4552 4870 4566 4922
rect 4590 4870 4604 4922
rect 4604 4870 4616 4922
rect 4616 4870 4646 4922
rect 4670 4870 4680 4922
rect 4680 4870 4726 4922
rect 4430 4868 4486 4870
rect 4510 4868 4566 4870
rect 4590 4868 4646 4870
rect 4670 4868 4726 4870
rect 4430 3834 4486 3836
rect 4510 3834 4566 3836
rect 4590 3834 4646 3836
rect 4670 3834 4726 3836
rect 4430 3782 4476 3834
rect 4476 3782 4486 3834
rect 4510 3782 4540 3834
rect 4540 3782 4552 3834
rect 4552 3782 4566 3834
rect 4590 3782 4604 3834
rect 4604 3782 4616 3834
rect 4616 3782 4646 3834
rect 4670 3782 4680 3834
rect 4680 3782 4726 3834
rect 4430 3780 4486 3782
rect 4510 3780 4566 3782
rect 4590 3780 4646 3782
rect 4670 3780 4726 3782
rect 4430 2746 4486 2748
rect 4510 2746 4566 2748
rect 4590 2746 4646 2748
rect 4670 2746 4726 2748
rect 4430 2694 4476 2746
rect 4476 2694 4486 2746
rect 4510 2694 4540 2746
rect 4540 2694 4552 2746
rect 4552 2694 4566 2746
rect 4590 2694 4604 2746
rect 4604 2694 4616 2746
rect 4616 2694 4646 2746
rect 4670 2694 4680 2746
rect 4680 2694 4726 2746
rect 4430 2692 4486 2694
rect 4510 2692 4566 2694
rect 4590 2692 4646 2694
rect 4670 2692 4726 2694
rect 7904 13082 7960 13084
rect 7984 13082 8040 13084
rect 8064 13082 8120 13084
rect 8144 13082 8200 13084
rect 7904 13030 7950 13082
rect 7950 13030 7960 13082
rect 7984 13030 8014 13082
rect 8014 13030 8026 13082
rect 8026 13030 8040 13082
rect 8064 13030 8078 13082
rect 8078 13030 8090 13082
rect 8090 13030 8120 13082
rect 8144 13030 8154 13082
rect 8154 13030 8200 13082
rect 7904 13028 7960 13030
rect 7984 13028 8040 13030
rect 8064 13028 8120 13030
rect 8144 13028 8200 13030
rect 7904 11994 7960 11996
rect 7984 11994 8040 11996
rect 8064 11994 8120 11996
rect 8144 11994 8200 11996
rect 7904 11942 7950 11994
rect 7950 11942 7960 11994
rect 7984 11942 8014 11994
rect 8014 11942 8026 11994
rect 8026 11942 8040 11994
rect 8064 11942 8078 11994
rect 8078 11942 8090 11994
rect 8090 11942 8120 11994
rect 8144 11942 8154 11994
rect 8154 11942 8200 11994
rect 7904 11940 7960 11942
rect 7984 11940 8040 11942
rect 8064 11940 8120 11942
rect 8144 11940 8200 11942
rect 7904 10906 7960 10908
rect 7984 10906 8040 10908
rect 8064 10906 8120 10908
rect 8144 10906 8200 10908
rect 7904 10854 7950 10906
rect 7950 10854 7960 10906
rect 7984 10854 8014 10906
rect 8014 10854 8026 10906
rect 8026 10854 8040 10906
rect 8064 10854 8078 10906
rect 8078 10854 8090 10906
rect 8090 10854 8120 10906
rect 8144 10854 8154 10906
rect 8154 10854 8200 10906
rect 7904 10852 7960 10854
rect 7984 10852 8040 10854
rect 8064 10852 8120 10854
rect 8144 10852 8200 10854
rect 7904 9818 7960 9820
rect 7984 9818 8040 9820
rect 8064 9818 8120 9820
rect 8144 9818 8200 9820
rect 7904 9766 7950 9818
rect 7950 9766 7960 9818
rect 7984 9766 8014 9818
rect 8014 9766 8026 9818
rect 8026 9766 8040 9818
rect 8064 9766 8078 9818
rect 8078 9766 8090 9818
rect 8090 9766 8120 9818
rect 8144 9766 8154 9818
rect 8154 9766 8200 9818
rect 7904 9764 7960 9766
rect 7984 9764 8040 9766
rect 8064 9764 8120 9766
rect 8144 9764 8200 9766
rect 11378 15802 11434 15804
rect 11458 15802 11514 15804
rect 11538 15802 11594 15804
rect 11618 15802 11674 15804
rect 11378 15750 11424 15802
rect 11424 15750 11434 15802
rect 11458 15750 11488 15802
rect 11488 15750 11500 15802
rect 11500 15750 11514 15802
rect 11538 15750 11552 15802
rect 11552 15750 11564 15802
rect 11564 15750 11594 15802
rect 11618 15750 11628 15802
rect 11628 15750 11674 15802
rect 11378 15748 11434 15750
rect 11458 15748 11514 15750
rect 11538 15748 11594 15750
rect 11618 15748 11674 15750
rect 14852 16346 14908 16348
rect 14932 16346 14988 16348
rect 15012 16346 15068 16348
rect 15092 16346 15148 16348
rect 14852 16294 14898 16346
rect 14898 16294 14908 16346
rect 14932 16294 14962 16346
rect 14962 16294 14974 16346
rect 14974 16294 14988 16346
rect 15012 16294 15026 16346
rect 15026 16294 15038 16346
rect 15038 16294 15068 16346
rect 15092 16294 15102 16346
rect 15102 16294 15148 16346
rect 14852 16292 14908 16294
rect 14932 16292 14988 16294
rect 15012 16292 15068 16294
rect 15092 16292 15148 16294
rect 7904 8730 7960 8732
rect 7984 8730 8040 8732
rect 8064 8730 8120 8732
rect 8144 8730 8200 8732
rect 7904 8678 7950 8730
rect 7950 8678 7960 8730
rect 7984 8678 8014 8730
rect 8014 8678 8026 8730
rect 8026 8678 8040 8730
rect 8064 8678 8078 8730
rect 8078 8678 8090 8730
rect 8090 8678 8120 8730
rect 8144 8678 8154 8730
rect 8154 8678 8200 8730
rect 7904 8676 7960 8678
rect 7984 8676 8040 8678
rect 8064 8676 8120 8678
rect 8144 8676 8200 8678
rect 11378 14714 11434 14716
rect 11458 14714 11514 14716
rect 11538 14714 11594 14716
rect 11618 14714 11674 14716
rect 11378 14662 11424 14714
rect 11424 14662 11434 14714
rect 11458 14662 11488 14714
rect 11488 14662 11500 14714
rect 11500 14662 11514 14714
rect 11538 14662 11552 14714
rect 11552 14662 11564 14714
rect 11564 14662 11594 14714
rect 11618 14662 11628 14714
rect 11628 14662 11674 14714
rect 11378 14660 11434 14662
rect 11458 14660 11514 14662
rect 11538 14660 11594 14662
rect 11618 14660 11674 14662
rect 11378 13626 11434 13628
rect 11458 13626 11514 13628
rect 11538 13626 11594 13628
rect 11618 13626 11674 13628
rect 11378 13574 11424 13626
rect 11424 13574 11434 13626
rect 11458 13574 11488 13626
rect 11488 13574 11500 13626
rect 11500 13574 11514 13626
rect 11538 13574 11552 13626
rect 11552 13574 11564 13626
rect 11564 13574 11594 13626
rect 11618 13574 11628 13626
rect 11628 13574 11674 13626
rect 11378 13572 11434 13574
rect 11458 13572 11514 13574
rect 11538 13572 11594 13574
rect 11618 13572 11674 13574
rect 11150 13232 11206 13288
rect 11378 12538 11434 12540
rect 11458 12538 11514 12540
rect 11538 12538 11594 12540
rect 11618 12538 11674 12540
rect 11378 12486 11424 12538
rect 11424 12486 11434 12538
rect 11458 12486 11488 12538
rect 11488 12486 11500 12538
rect 11500 12486 11514 12538
rect 11538 12486 11552 12538
rect 11552 12486 11564 12538
rect 11564 12486 11594 12538
rect 11618 12486 11628 12538
rect 11628 12486 11674 12538
rect 11378 12484 11434 12486
rect 11458 12484 11514 12486
rect 11538 12484 11594 12486
rect 11618 12484 11674 12486
rect 11378 11450 11434 11452
rect 11458 11450 11514 11452
rect 11538 11450 11594 11452
rect 11618 11450 11674 11452
rect 11378 11398 11424 11450
rect 11424 11398 11434 11450
rect 11458 11398 11488 11450
rect 11488 11398 11500 11450
rect 11500 11398 11514 11450
rect 11538 11398 11552 11450
rect 11552 11398 11564 11450
rect 11564 11398 11594 11450
rect 11618 11398 11628 11450
rect 11628 11398 11674 11450
rect 11378 11396 11434 11398
rect 11458 11396 11514 11398
rect 11538 11396 11594 11398
rect 11618 11396 11674 11398
rect 11378 10362 11434 10364
rect 11458 10362 11514 10364
rect 11538 10362 11594 10364
rect 11618 10362 11674 10364
rect 11378 10310 11424 10362
rect 11424 10310 11434 10362
rect 11458 10310 11488 10362
rect 11488 10310 11500 10362
rect 11500 10310 11514 10362
rect 11538 10310 11552 10362
rect 11552 10310 11564 10362
rect 11564 10310 11594 10362
rect 11618 10310 11628 10362
rect 11628 10310 11674 10362
rect 11378 10308 11434 10310
rect 11458 10308 11514 10310
rect 11538 10308 11594 10310
rect 11618 10308 11674 10310
rect 11378 9274 11434 9276
rect 11458 9274 11514 9276
rect 11538 9274 11594 9276
rect 11618 9274 11674 9276
rect 11378 9222 11424 9274
rect 11424 9222 11434 9274
rect 11458 9222 11488 9274
rect 11488 9222 11500 9274
rect 11500 9222 11514 9274
rect 11538 9222 11552 9274
rect 11552 9222 11564 9274
rect 11564 9222 11594 9274
rect 11618 9222 11628 9274
rect 11628 9222 11674 9274
rect 11378 9220 11434 9222
rect 11458 9220 11514 9222
rect 11538 9220 11594 9222
rect 11618 9220 11674 9222
rect 7904 7642 7960 7644
rect 7984 7642 8040 7644
rect 8064 7642 8120 7644
rect 8144 7642 8200 7644
rect 7904 7590 7950 7642
rect 7950 7590 7960 7642
rect 7984 7590 8014 7642
rect 8014 7590 8026 7642
rect 8026 7590 8040 7642
rect 8064 7590 8078 7642
rect 8078 7590 8090 7642
rect 8090 7590 8120 7642
rect 8144 7590 8154 7642
rect 8154 7590 8200 7642
rect 7904 7588 7960 7590
rect 7984 7588 8040 7590
rect 8064 7588 8120 7590
rect 8144 7588 8200 7590
rect 11378 8186 11434 8188
rect 11458 8186 11514 8188
rect 11538 8186 11594 8188
rect 11618 8186 11674 8188
rect 11378 8134 11424 8186
rect 11424 8134 11434 8186
rect 11458 8134 11488 8186
rect 11488 8134 11500 8186
rect 11500 8134 11514 8186
rect 11538 8134 11552 8186
rect 11552 8134 11564 8186
rect 11564 8134 11594 8186
rect 11618 8134 11628 8186
rect 11628 8134 11674 8186
rect 11378 8132 11434 8134
rect 11458 8132 11514 8134
rect 11538 8132 11594 8134
rect 11618 8132 11674 8134
rect 11378 7098 11434 7100
rect 11458 7098 11514 7100
rect 11538 7098 11594 7100
rect 11618 7098 11674 7100
rect 11378 7046 11424 7098
rect 11424 7046 11434 7098
rect 11458 7046 11488 7098
rect 11488 7046 11500 7098
rect 11500 7046 11514 7098
rect 11538 7046 11552 7098
rect 11552 7046 11564 7098
rect 11564 7046 11594 7098
rect 11618 7046 11628 7098
rect 11628 7046 11674 7098
rect 11378 7044 11434 7046
rect 11458 7044 11514 7046
rect 11538 7044 11594 7046
rect 11618 7044 11674 7046
rect 7746 6704 7802 6760
rect 7904 6554 7960 6556
rect 7984 6554 8040 6556
rect 8064 6554 8120 6556
rect 8144 6554 8200 6556
rect 7904 6502 7950 6554
rect 7950 6502 7960 6554
rect 7984 6502 8014 6554
rect 8014 6502 8026 6554
rect 8026 6502 8040 6554
rect 8064 6502 8078 6554
rect 8078 6502 8090 6554
rect 8090 6502 8120 6554
rect 8144 6502 8154 6554
rect 8154 6502 8200 6554
rect 7904 6500 7960 6502
rect 7984 6500 8040 6502
rect 8064 6500 8120 6502
rect 8144 6500 8200 6502
rect 14094 6840 14150 6896
rect 11378 6010 11434 6012
rect 11458 6010 11514 6012
rect 11538 6010 11594 6012
rect 11618 6010 11674 6012
rect 11378 5958 11424 6010
rect 11424 5958 11434 6010
rect 11458 5958 11488 6010
rect 11488 5958 11500 6010
rect 11500 5958 11514 6010
rect 11538 5958 11552 6010
rect 11552 5958 11564 6010
rect 11564 5958 11594 6010
rect 11618 5958 11628 6010
rect 11628 5958 11674 6010
rect 11378 5956 11434 5958
rect 11458 5956 11514 5958
rect 11538 5956 11594 5958
rect 11618 5956 11674 5958
rect 7904 5466 7960 5468
rect 7984 5466 8040 5468
rect 8064 5466 8120 5468
rect 8144 5466 8200 5468
rect 7904 5414 7950 5466
rect 7950 5414 7960 5466
rect 7984 5414 8014 5466
rect 8014 5414 8026 5466
rect 8026 5414 8040 5466
rect 8064 5414 8078 5466
rect 8078 5414 8090 5466
rect 8090 5414 8120 5466
rect 8144 5414 8154 5466
rect 8154 5414 8200 5466
rect 7904 5412 7960 5414
rect 7984 5412 8040 5414
rect 8064 5412 8120 5414
rect 8144 5412 8200 5414
rect 11378 4922 11434 4924
rect 11458 4922 11514 4924
rect 11538 4922 11594 4924
rect 11618 4922 11674 4924
rect 11378 4870 11424 4922
rect 11424 4870 11434 4922
rect 11458 4870 11488 4922
rect 11488 4870 11500 4922
rect 11500 4870 11514 4922
rect 11538 4870 11552 4922
rect 11552 4870 11564 4922
rect 11564 4870 11594 4922
rect 11618 4870 11628 4922
rect 11628 4870 11674 4922
rect 11378 4868 11434 4870
rect 11458 4868 11514 4870
rect 11538 4868 11594 4870
rect 11618 4868 11674 4870
rect 7904 4378 7960 4380
rect 7984 4378 8040 4380
rect 8064 4378 8120 4380
rect 8144 4378 8200 4380
rect 7904 4326 7950 4378
rect 7950 4326 7960 4378
rect 7984 4326 8014 4378
rect 8014 4326 8026 4378
rect 8026 4326 8040 4378
rect 8064 4326 8078 4378
rect 8078 4326 8090 4378
rect 8090 4326 8120 4378
rect 8144 4326 8154 4378
rect 8154 4326 8200 4378
rect 7904 4324 7960 4326
rect 7984 4324 8040 4326
rect 8064 4324 8120 4326
rect 8144 4324 8200 4326
rect 7904 3290 7960 3292
rect 7984 3290 8040 3292
rect 8064 3290 8120 3292
rect 8144 3290 8200 3292
rect 7904 3238 7950 3290
rect 7950 3238 7960 3290
rect 7984 3238 8014 3290
rect 8014 3238 8026 3290
rect 8026 3238 8040 3290
rect 8064 3238 8078 3290
rect 8078 3238 8090 3290
rect 8090 3238 8120 3290
rect 8144 3238 8154 3290
rect 8154 3238 8200 3290
rect 7904 3236 7960 3238
rect 7984 3236 8040 3238
rect 8064 3236 8120 3238
rect 8144 3236 8200 3238
rect 11378 3834 11434 3836
rect 11458 3834 11514 3836
rect 11538 3834 11594 3836
rect 11618 3834 11674 3836
rect 11378 3782 11424 3834
rect 11424 3782 11434 3834
rect 11458 3782 11488 3834
rect 11488 3782 11500 3834
rect 11500 3782 11514 3834
rect 11538 3782 11552 3834
rect 11552 3782 11564 3834
rect 11564 3782 11594 3834
rect 11618 3782 11628 3834
rect 11628 3782 11674 3834
rect 11378 3780 11434 3782
rect 11458 3780 11514 3782
rect 11538 3780 11594 3782
rect 11618 3780 11674 3782
rect 14852 15258 14908 15260
rect 14932 15258 14988 15260
rect 15012 15258 15068 15260
rect 15092 15258 15148 15260
rect 14852 15206 14898 15258
rect 14898 15206 14908 15258
rect 14932 15206 14962 15258
rect 14962 15206 14974 15258
rect 14974 15206 14988 15258
rect 15012 15206 15026 15258
rect 15026 15206 15038 15258
rect 15038 15206 15068 15258
rect 15092 15206 15102 15258
rect 15102 15206 15148 15258
rect 14852 15204 14908 15206
rect 14932 15204 14988 15206
rect 15012 15204 15068 15206
rect 15092 15204 15148 15206
rect 14852 14170 14908 14172
rect 14932 14170 14988 14172
rect 15012 14170 15068 14172
rect 15092 14170 15148 14172
rect 14852 14118 14898 14170
rect 14898 14118 14908 14170
rect 14932 14118 14962 14170
rect 14962 14118 14974 14170
rect 14974 14118 14988 14170
rect 15012 14118 15026 14170
rect 15026 14118 15038 14170
rect 15038 14118 15068 14170
rect 15092 14118 15102 14170
rect 15102 14118 15148 14170
rect 14852 14116 14908 14118
rect 14932 14116 14988 14118
rect 15012 14116 15068 14118
rect 15092 14116 15148 14118
rect 14852 13082 14908 13084
rect 14932 13082 14988 13084
rect 15012 13082 15068 13084
rect 15092 13082 15148 13084
rect 14852 13030 14898 13082
rect 14898 13030 14908 13082
rect 14932 13030 14962 13082
rect 14962 13030 14974 13082
rect 14974 13030 14988 13082
rect 15012 13030 15026 13082
rect 15026 13030 15038 13082
rect 15038 13030 15068 13082
rect 15092 13030 15102 13082
rect 15102 13030 15148 13082
rect 14852 13028 14908 13030
rect 14932 13028 14988 13030
rect 15012 13028 15068 13030
rect 15092 13028 15148 13030
rect 14852 11994 14908 11996
rect 14932 11994 14988 11996
rect 15012 11994 15068 11996
rect 15092 11994 15148 11996
rect 14852 11942 14898 11994
rect 14898 11942 14908 11994
rect 14932 11942 14962 11994
rect 14962 11942 14974 11994
rect 14974 11942 14988 11994
rect 15012 11942 15026 11994
rect 15026 11942 15038 11994
rect 15038 11942 15068 11994
rect 15092 11942 15102 11994
rect 15102 11942 15148 11994
rect 14852 11940 14908 11942
rect 14932 11940 14988 11942
rect 15012 11940 15068 11942
rect 15092 11940 15148 11942
rect 14852 10906 14908 10908
rect 14932 10906 14988 10908
rect 15012 10906 15068 10908
rect 15092 10906 15148 10908
rect 14852 10854 14898 10906
rect 14898 10854 14908 10906
rect 14932 10854 14962 10906
rect 14962 10854 14974 10906
rect 14974 10854 14988 10906
rect 15012 10854 15026 10906
rect 15026 10854 15038 10906
rect 15038 10854 15068 10906
rect 15092 10854 15102 10906
rect 15102 10854 15148 10906
rect 14852 10852 14908 10854
rect 14932 10852 14988 10854
rect 15012 10852 15068 10854
rect 15092 10852 15148 10854
rect 14852 9818 14908 9820
rect 14932 9818 14988 9820
rect 15012 9818 15068 9820
rect 15092 9818 15148 9820
rect 14852 9766 14898 9818
rect 14898 9766 14908 9818
rect 14932 9766 14962 9818
rect 14962 9766 14974 9818
rect 14974 9766 14988 9818
rect 15012 9766 15026 9818
rect 15026 9766 15038 9818
rect 15038 9766 15068 9818
rect 15092 9766 15102 9818
rect 15102 9766 15148 9818
rect 14852 9764 14908 9766
rect 14932 9764 14988 9766
rect 15012 9764 15068 9766
rect 15092 9764 15148 9766
rect 14852 8730 14908 8732
rect 14932 8730 14988 8732
rect 15012 8730 15068 8732
rect 15092 8730 15148 8732
rect 14852 8678 14898 8730
rect 14898 8678 14908 8730
rect 14932 8678 14962 8730
rect 14962 8678 14974 8730
rect 14974 8678 14988 8730
rect 15012 8678 15026 8730
rect 15026 8678 15038 8730
rect 15038 8678 15068 8730
rect 15092 8678 15102 8730
rect 15102 8678 15148 8730
rect 14852 8676 14908 8678
rect 14932 8676 14988 8678
rect 15012 8676 15068 8678
rect 15092 8676 15148 8678
rect 14852 7642 14908 7644
rect 14932 7642 14988 7644
rect 15012 7642 15068 7644
rect 15092 7642 15148 7644
rect 14852 7590 14898 7642
rect 14898 7590 14908 7642
rect 14932 7590 14962 7642
rect 14962 7590 14974 7642
rect 14974 7590 14988 7642
rect 15012 7590 15026 7642
rect 15026 7590 15038 7642
rect 15038 7590 15068 7642
rect 15092 7590 15102 7642
rect 15102 7590 15148 7642
rect 14852 7588 14908 7590
rect 14932 7588 14988 7590
rect 15012 7588 15068 7590
rect 15092 7588 15148 7590
rect 21800 27226 21856 27228
rect 21880 27226 21936 27228
rect 21960 27226 22016 27228
rect 22040 27226 22096 27228
rect 21800 27174 21846 27226
rect 21846 27174 21856 27226
rect 21880 27174 21910 27226
rect 21910 27174 21922 27226
rect 21922 27174 21936 27226
rect 21960 27174 21974 27226
rect 21974 27174 21986 27226
rect 21986 27174 22016 27226
rect 22040 27174 22050 27226
rect 22050 27174 22096 27226
rect 21800 27172 21856 27174
rect 21880 27172 21936 27174
rect 21960 27172 22016 27174
rect 22040 27172 22096 27174
rect 18326 26682 18382 26684
rect 18406 26682 18462 26684
rect 18486 26682 18542 26684
rect 18566 26682 18622 26684
rect 18326 26630 18372 26682
rect 18372 26630 18382 26682
rect 18406 26630 18436 26682
rect 18436 26630 18448 26682
rect 18448 26630 18462 26682
rect 18486 26630 18500 26682
rect 18500 26630 18512 26682
rect 18512 26630 18542 26682
rect 18566 26630 18576 26682
rect 18576 26630 18622 26682
rect 18326 26628 18382 26630
rect 18406 26628 18462 26630
rect 18486 26628 18542 26630
rect 18566 26628 18622 26630
rect 25274 26682 25330 26684
rect 25354 26682 25410 26684
rect 25434 26682 25490 26684
rect 25514 26682 25570 26684
rect 25274 26630 25320 26682
rect 25320 26630 25330 26682
rect 25354 26630 25384 26682
rect 25384 26630 25396 26682
rect 25396 26630 25410 26682
rect 25434 26630 25448 26682
rect 25448 26630 25460 26682
rect 25460 26630 25490 26682
rect 25514 26630 25524 26682
rect 25524 26630 25570 26682
rect 25274 26628 25330 26630
rect 25354 26628 25410 26630
rect 25434 26628 25490 26630
rect 25514 26628 25570 26630
rect 21800 26138 21856 26140
rect 21880 26138 21936 26140
rect 21960 26138 22016 26140
rect 22040 26138 22096 26140
rect 21800 26086 21846 26138
rect 21846 26086 21856 26138
rect 21880 26086 21910 26138
rect 21910 26086 21922 26138
rect 21922 26086 21936 26138
rect 21960 26086 21974 26138
rect 21974 26086 21986 26138
rect 21986 26086 22016 26138
rect 22040 26086 22050 26138
rect 22050 26086 22096 26138
rect 21800 26084 21856 26086
rect 21880 26084 21936 26086
rect 21960 26084 22016 26086
rect 22040 26084 22096 26086
rect 18326 25594 18382 25596
rect 18406 25594 18462 25596
rect 18486 25594 18542 25596
rect 18566 25594 18622 25596
rect 18326 25542 18372 25594
rect 18372 25542 18382 25594
rect 18406 25542 18436 25594
rect 18436 25542 18448 25594
rect 18448 25542 18462 25594
rect 18486 25542 18500 25594
rect 18500 25542 18512 25594
rect 18512 25542 18542 25594
rect 18566 25542 18576 25594
rect 18576 25542 18622 25594
rect 18326 25540 18382 25542
rect 18406 25540 18462 25542
rect 18486 25540 18542 25542
rect 18566 25540 18622 25542
rect 25274 25594 25330 25596
rect 25354 25594 25410 25596
rect 25434 25594 25490 25596
rect 25514 25594 25570 25596
rect 25274 25542 25320 25594
rect 25320 25542 25330 25594
rect 25354 25542 25384 25594
rect 25384 25542 25396 25594
rect 25396 25542 25410 25594
rect 25434 25542 25448 25594
rect 25448 25542 25460 25594
rect 25460 25542 25490 25594
rect 25514 25542 25524 25594
rect 25524 25542 25570 25594
rect 25274 25540 25330 25542
rect 25354 25540 25410 25542
rect 25434 25540 25490 25542
rect 25514 25540 25570 25542
rect 21800 25050 21856 25052
rect 21880 25050 21936 25052
rect 21960 25050 22016 25052
rect 22040 25050 22096 25052
rect 21800 24998 21846 25050
rect 21846 24998 21856 25050
rect 21880 24998 21910 25050
rect 21910 24998 21922 25050
rect 21922 24998 21936 25050
rect 21960 24998 21974 25050
rect 21974 24998 21986 25050
rect 21986 24998 22016 25050
rect 22040 24998 22050 25050
rect 22050 24998 22096 25050
rect 21800 24996 21856 24998
rect 21880 24996 21936 24998
rect 21960 24996 22016 24998
rect 22040 24996 22096 24998
rect 18326 24506 18382 24508
rect 18406 24506 18462 24508
rect 18486 24506 18542 24508
rect 18566 24506 18622 24508
rect 18326 24454 18372 24506
rect 18372 24454 18382 24506
rect 18406 24454 18436 24506
rect 18436 24454 18448 24506
rect 18448 24454 18462 24506
rect 18486 24454 18500 24506
rect 18500 24454 18512 24506
rect 18512 24454 18542 24506
rect 18566 24454 18576 24506
rect 18576 24454 18622 24506
rect 18326 24452 18382 24454
rect 18406 24452 18462 24454
rect 18486 24452 18542 24454
rect 18566 24452 18622 24454
rect 25274 24506 25330 24508
rect 25354 24506 25410 24508
rect 25434 24506 25490 24508
rect 25514 24506 25570 24508
rect 25274 24454 25320 24506
rect 25320 24454 25330 24506
rect 25354 24454 25384 24506
rect 25384 24454 25396 24506
rect 25396 24454 25410 24506
rect 25434 24454 25448 24506
rect 25448 24454 25460 24506
rect 25460 24454 25490 24506
rect 25514 24454 25524 24506
rect 25524 24454 25570 24506
rect 25274 24452 25330 24454
rect 25354 24452 25410 24454
rect 25434 24452 25490 24454
rect 25514 24452 25570 24454
rect 21800 23962 21856 23964
rect 21880 23962 21936 23964
rect 21960 23962 22016 23964
rect 22040 23962 22096 23964
rect 21800 23910 21846 23962
rect 21846 23910 21856 23962
rect 21880 23910 21910 23962
rect 21910 23910 21922 23962
rect 21922 23910 21936 23962
rect 21960 23910 21974 23962
rect 21974 23910 21986 23962
rect 21986 23910 22016 23962
rect 22040 23910 22050 23962
rect 22050 23910 22096 23962
rect 21800 23908 21856 23910
rect 21880 23908 21936 23910
rect 21960 23908 22016 23910
rect 22040 23908 22096 23910
rect 18326 23418 18382 23420
rect 18406 23418 18462 23420
rect 18486 23418 18542 23420
rect 18566 23418 18622 23420
rect 18326 23366 18372 23418
rect 18372 23366 18382 23418
rect 18406 23366 18436 23418
rect 18436 23366 18448 23418
rect 18448 23366 18462 23418
rect 18486 23366 18500 23418
rect 18500 23366 18512 23418
rect 18512 23366 18542 23418
rect 18566 23366 18576 23418
rect 18576 23366 18622 23418
rect 18326 23364 18382 23366
rect 18406 23364 18462 23366
rect 18486 23364 18542 23366
rect 18566 23364 18622 23366
rect 25274 23418 25330 23420
rect 25354 23418 25410 23420
rect 25434 23418 25490 23420
rect 25514 23418 25570 23420
rect 25274 23366 25320 23418
rect 25320 23366 25330 23418
rect 25354 23366 25384 23418
rect 25384 23366 25396 23418
rect 25396 23366 25410 23418
rect 25434 23366 25448 23418
rect 25448 23366 25460 23418
rect 25460 23366 25490 23418
rect 25514 23366 25524 23418
rect 25524 23366 25570 23418
rect 25274 23364 25330 23366
rect 25354 23364 25410 23366
rect 25434 23364 25490 23366
rect 25514 23364 25570 23366
rect 21800 22874 21856 22876
rect 21880 22874 21936 22876
rect 21960 22874 22016 22876
rect 22040 22874 22096 22876
rect 21800 22822 21846 22874
rect 21846 22822 21856 22874
rect 21880 22822 21910 22874
rect 21910 22822 21922 22874
rect 21922 22822 21936 22874
rect 21960 22822 21974 22874
rect 21974 22822 21986 22874
rect 21986 22822 22016 22874
rect 22040 22822 22050 22874
rect 22050 22822 22096 22874
rect 21800 22820 21856 22822
rect 21880 22820 21936 22822
rect 21960 22820 22016 22822
rect 22040 22820 22096 22822
rect 18326 22330 18382 22332
rect 18406 22330 18462 22332
rect 18486 22330 18542 22332
rect 18566 22330 18622 22332
rect 18326 22278 18372 22330
rect 18372 22278 18382 22330
rect 18406 22278 18436 22330
rect 18436 22278 18448 22330
rect 18448 22278 18462 22330
rect 18486 22278 18500 22330
rect 18500 22278 18512 22330
rect 18512 22278 18542 22330
rect 18566 22278 18576 22330
rect 18576 22278 18622 22330
rect 18326 22276 18382 22278
rect 18406 22276 18462 22278
rect 18486 22276 18542 22278
rect 18566 22276 18622 22278
rect 25274 22330 25330 22332
rect 25354 22330 25410 22332
rect 25434 22330 25490 22332
rect 25514 22330 25570 22332
rect 25274 22278 25320 22330
rect 25320 22278 25330 22330
rect 25354 22278 25384 22330
rect 25384 22278 25396 22330
rect 25396 22278 25410 22330
rect 25434 22278 25448 22330
rect 25448 22278 25460 22330
rect 25460 22278 25490 22330
rect 25514 22278 25524 22330
rect 25524 22278 25570 22330
rect 25274 22276 25330 22278
rect 25354 22276 25410 22278
rect 25434 22276 25490 22278
rect 25514 22276 25570 22278
rect 21800 21786 21856 21788
rect 21880 21786 21936 21788
rect 21960 21786 22016 21788
rect 22040 21786 22096 21788
rect 21800 21734 21846 21786
rect 21846 21734 21856 21786
rect 21880 21734 21910 21786
rect 21910 21734 21922 21786
rect 21922 21734 21936 21786
rect 21960 21734 21974 21786
rect 21974 21734 21986 21786
rect 21986 21734 22016 21786
rect 22040 21734 22050 21786
rect 22050 21734 22096 21786
rect 21800 21732 21856 21734
rect 21880 21732 21936 21734
rect 21960 21732 22016 21734
rect 22040 21732 22096 21734
rect 18326 21242 18382 21244
rect 18406 21242 18462 21244
rect 18486 21242 18542 21244
rect 18566 21242 18622 21244
rect 18326 21190 18372 21242
rect 18372 21190 18382 21242
rect 18406 21190 18436 21242
rect 18436 21190 18448 21242
rect 18448 21190 18462 21242
rect 18486 21190 18500 21242
rect 18500 21190 18512 21242
rect 18512 21190 18542 21242
rect 18566 21190 18576 21242
rect 18576 21190 18622 21242
rect 18326 21188 18382 21190
rect 18406 21188 18462 21190
rect 18486 21188 18542 21190
rect 18566 21188 18622 21190
rect 25274 21242 25330 21244
rect 25354 21242 25410 21244
rect 25434 21242 25490 21244
rect 25514 21242 25570 21244
rect 25274 21190 25320 21242
rect 25320 21190 25330 21242
rect 25354 21190 25384 21242
rect 25384 21190 25396 21242
rect 25396 21190 25410 21242
rect 25434 21190 25448 21242
rect 25448 21190 25460 21242
rect 25460 21190 25490 21242
rect 25514 21190 25524 21242
rect 25524 21190 25570 21242
rect 25274 21188 25330 21190
rect 25354 21188 25410 21190
rect 25434 21188 25490 21190
rect 25514 21188 25570 21190
rect 21800 20698 21856 20700
rect 21880 20698 21936 20700
rect 21960 20698 22016 20700
rect 22040 20698 22096 20700
rect 21800 20646 21846 20698
rect 21846 20646 21856 20698
rect 21880 20646 21910 20698
rect 21910 20646 21922 20698
rect 21922 20646 21936 20698
rect 21960 20646 21974 20698
rect 21974 20646 21986 20698
rect 21986 20646 22016 20698
rect 22040 20646 22050 20698
rect 22050 20646 22096 20698
rect 21800 20644 21856 20646
rect 21880 20644 21936 20646
rect 21960 20644 22016 20646
rect 22040 20644 22096 20646
rect 18326 20154 18382 20156
rect 18406 20154 18462 20156
rect 18486 20154 18542 20156
rect 18566 20154 18622 20156
rect 18326 20102 18372 20154
rect 18372 20102 18382 20154
rect 18406 20102 18436 20154
rect 18436 20102 18448 20154
rect 18448 20102 18462 20154
rect 18486 20102 18500 20154
rect 18500 20102 18512 20154
rect 18512 20102 18542 20154
rect 18566 20102 18576 20154
rect 18576 20102 18622 20154
rect 18326 20100 18382 20102
rect 18406 20100 18462 20102
rect 18486 20100 18542 20102
rect 18566 20100 18622 20102
rect 25274 20154 25330 20156
rect 25354 20154 25410 20156
rect 25434 20154 25490 20156
rect 25514 20154 25570 20156
rect 25274 20102 25320 20154
rect 25320 20102 25330 20154
rect 25354 20102 25384 20154
rect 25384 20102 25396 20154
rect 25396 20102 25410 20154
rect 25434 20102 25448 20154
rect 25448 20102 25460 20154
rect 25460 20102 25490 20154
rect 25514 20102 25524 20154
rect 25524 20102 25570 20154
rect 25274 20100 25330 20102
rect 25354 20100 25410 20102
rect 25434 20100 25490 20102
rect 25514 20100 25570 20102
rect 21800 19610 21856 19612
rect 21880 19610 21936 19612
rect 21960 19610 22016 19612
rect 22040 19610 22096 19612
rect 21800 19558 21846 19610
rect 21846 19558 21856 19610
rect 21880 19558 21910 19610
rect 21910 19558 21922 19610
rect 21922 19558 21936 19610
rect 21960 19558 21974 19610
rect 21974 19558 21986 19610
rect 21986 19558 22016 19610
rect 22040 19558 22050 19610
rect 22050 19558 22096 19610
rect 21800 19556 21856 19558
rect 21880 19556 21936 19558
rect 21960 19556 22016 19558
rect 22040 19556 22096 19558
rect 18326 19066 18382 19068
rect 18406 19066 18462 19068
rect 18486 19066 18542 19068
rect 18566 19066 18622 19068
rect 18326 19014 18372 19066
rect 18372 19014 18382 19066
rect 18406 19014 18436 19066
rect 18436 19014 18448 19066
rect 18448 19014 18462 19066
rect 18486 19014 18500 19066
rect 18500 19014 18512 19066
rect 18512 19014 18542 19066
rect 18566 19014 18576 19066
rect 18576 19014 18622 19066
rect 18326 19012 18382 19014
rect 18406 19012 18462 19014
rect 18486 19012 18542 19014
rect 18566 19012 18622 19014
rect 25274 19066 25330 19068
rect 25354 19066 25410 19068
rect 25434 19066 25490 19068
rect 25514 19066 25570 19068
rect 25274 19014 25320 19066
rect 25320 19014 25330 19066
rect 25354 19014 25384 19066
rect 25384 19014 25396 19066
rect 25396 19014 25410 19066
rect 25434 19014 25448 19066
rect 25448 19014 25460 19066
rect 25460 19014 25490 19066
rect 25514 19014 25524 19066
rect 25524 19014 25570 19066
rect 25274 19012 25330 19014
rect 25354 19012 25410 19014
rect 25434 19012 25490 19014
rect 25514 19012 25570 19014
rect 21800 18522 21856 18524
rect 21880 18522 21936 18524
rect 21960 18522 22016 18524
rect 22040 18522 22096 18524
rect 21800 18470 21846 18522
rect 21846 18470 21856 18522
rect 21880 18470 21910 18522
rect 21910 18470 21922 18522
rect 21922 18470 21936 18522
rect 21960 18470 21974 18522
rect 21974 18470 21986 18522
rect 21986 18470 22016 18522
rect 22040 18470 22050 18522
rect 22050 18470 22096 18522
rect 21800 18468 21856 18470
rect 21880 18468 21936 18470
rect 21960 18468 22016 18470
rect 22040 18468 22096 18470
rect 18326 17978 18382 17980
rect 18406 17978 18462 17980
rect 18486 17978 18542 17980
rect 18566 17978 18622 17980
rect 18326 17926 18372 17978
rect 18372 17926 18382 17978
rect 18406 17926 18436 17978
rect 18436 17926 18448 17978
rect 18448 17926 18462 17978
rect 18486 17926 18500 17978
rect 18500 17926 18512 17978
rect 18512 17926 18542 17978
rect 18566 17926 18576 17978
rect 18576 17926 18622 17978
rect 18326 17924 18382 17926
rect 18406 17924 18462 17926
rect 18486 17924 18542 17926
rect 18566 17924 18622 17926
rect 25274 17978 25330 17980
rect 25354 17978 25410 17980
rect 25434 17978 25490 17980
rect 25514 17978 25570 17980
rect 25274 17926 25320 17978
rect 25320 17926 25330 17978
rect 25354 17926 25384 17978
rect 25384 17926 25396 17978
rect 25396 17926 25410 17978
rect 25434 17926 25448 17978
rect 25448 17926 25460 17978
rect 25460 17926 25490 17978
rect 25514 17926 25524 17978
rect 25524 17926 25570 17978
rect 25274 17924 25330 17926
rect 25354 17924 25410 17926
rect 25434 17924 25490 17926
rect 25514 17924 25570 17926
rect 21800 17434 21856 17436
rect 21880 17434 21936 17436
rect 21960 17434 22016 17436
rect 22040 17434 22096 17436
rect 21800 17382 21846 17434
rect 21846 17382 21856 17434
rect 21880 17382 21910 17434
rect 21910 17382 21922 17434
rect 21922 17382 21936 17434
rect 21960 17382 21974 17434
rect 21974 17382 21986 17434
rect 21986 17382 22016 17434
rect 22040 17382 22050 17434
rect 22050 17382 22096 17434
rect 21800 17380 21856 17382
rect 21880 17380 21936 17382
rect 21960 17380 22016 17382
rect 22040 17380 22096 17382
rect 28170 17040 28226 17096
rect 18326 16890 18382 16892
rect 18406 16890 18462 16892
rect 18486 16890 18542 16892
rect 18566 16890 18622 16892
rect 18326 16838 18372 16890
rect 18372 16838 18382 16890
rect 18406 16838 18436 16890
rect 18436 16838 18448 16890
rect 18448 16838 18462 16890
rect 18486 16838 18500 16890
rect 18500 16838 18512 16890
rect 18512 16838 18542 16890
rect 18566 16838 18576 16890
rect 18576 16838 18622 16890
rect 18326 16836 18382 16838
rect 18406 16836 18462 16838
rect 18486 16836 18542 16838
rect 18566 16836 18622 16838
rect 25274 16890 25330 16892
rect 25354 16890 25410 16892
rect 25434 16890 25490 16892
rect 25514 16890 25570 16892
rect 25274 16838 25320 16890
rect 25320 16838 25330 16890
rect 25354 16838 25384 16890
rect 25384 16838 25396 16890
rect 25396 16838 25410 16890
rect 25434 16838 25448 16890
rect 25448 16838 25460 16890
rect 25460 16838 25490 16890
rect 25514 16838 25524 16890
rect 25524 16838 25570 16890
rect 25274 16836 25330 16838
rect 25354 16836 25410 16838
rect 25434 16836 25490 16838
rect 25514 16836 25570 16838
rect 21800 16346 21856 16348
rect 21880 16346 21936 16348
rect 21960 16346 22016 16348
rect 22040 16346 22096 16348
rect 21800 16294 21846 16346
rect 21846 16294 21856 16346
rect 21880 16294 21910 16346
rect 21910 16294 21922 16346
rect 21922 16294 21936 16346
rect 21960 16294 21974 16346
rect 21974 16294 21986 16346
rect 21986 16294 22016 16346
rect 22040 16294 22050 16346
rect 22050 16294 22096 16346
rect 21800 16292 21856 16294
rect 21880 16292 21936 16294
rect 21960 16292 22016 16294
rect 22040 16292 22096 16294
rect 18326 15802 18382 15804
rect 18406 15802 18462 15804
rect 18486 15802 18542 15804
rect 18566 15802 18622 15804
rect 18326 15750 18372 15802
rect 18372 15750 18382 15802
rect 18406 15750 18436 15802
rect 18436 15750 18448 15802
rect 18448 15750 18462 15802
rect 18486 15750 18500 15802
rect 18500 15750 18512 15802
rect 18512 15750 18542 15802
rect 18566 15750 18576 15802
rect 18576 15750 18622 15802
rect 18326 15748 18382 15750
rect 18406 15748 18462 15750
rect 18486 15748 18542 15750
rect 18566 15748 18622 15750
rect 25274 15802 25330 15804
rect 25354 15802 25410 15804
rect 25434 15802 25490 15804
rect 25514 15802 25570 15804
rect 25274 15750 25320 15802
rect 25320 15750 25330 15802
rect 25354 15750 25384 15802
rect 25384 15750 25396 15802
rect 25396 15750 25410 15802
rect 25434 15750 25448 15802
rect 25448 15750 25460 15802
rect 25460 15750 25490 15802
rect 25514 15750 25524 15802
rect 25524 15750 25570 15802
rect 25274 15748 25330 15750
rect 25354 15748 25410 15750
rect 25434 15748 25490 15750
rect 25514 15748 25570 15750
rect 21800 15258 21856 15260
rect 21880 15258 21936 15260
rect 21960 15258 22016 15260
rect 22040 15258 22096 15260
rect 21800 15206 21846 15258
rect 21846 15206 21856 15258
rect 21880 15206 21910 15258
rect 21910 15206 21922 15258
rect 21922 15206 21936 15258
rect 21960 15206 21974 15258
rect 21974 15206 21986 15258
rect 21986 15206 22016 15258
rect 22040 15206 22050 15258
rect 22050 15206 22096 15258
rect 21800 15204 21856 15206
rect 21880 15204 21936 15206
rect 21960 15204 22016 15206
rect 22040 15204 22096 15206
rect 18326 14714 18382 14716
rect 18406 14714 18462 14716
rect 18486 14714 18542 14716
rect 18566 14714 18622 14716
rect 18326 14662 18372 14714
rect 18372 14662 18382 14714
rect 18406 14662 18436 14714
rect 18436 14662 18448 14714
rect 18448 14662 18462 14714
rect 18486 14662 18500 14714
rect 18500 14662 18512 14714
rect 18512 14662 18542 14714
rect 18566 14662 18576 14714
rect 18576 14662 18622 14714
rect 18326 14660 18382 14662
rect 18406 14660 18462 14662
rect 18486 14660 18542 14662
rect 18566 14660 18622 14662
rect 25274 14714 25330 14716
rect 25354 14714 25410 14716
rect 25434 14714 25490 14716
rect 25514 14714 25570 14716
rect 25274 14662 25320 14714
rect 25320 14662 25330 14714
rect 25354 14662 25384 14714
rect 25384 14662 25396 14714
rect 25396 14662 25410 14714
rect 25434 14662 25448 14714
rect 25448 14662 25460 14714
rect 25460 14662 25490 14714
rect 25514 14662 25524 14714
rect 25524 14662 25570 14714
rect 25274 14660 25330 14662
rect 25354 14660 25410 14662
rect 25434 14660 25490 14662
rect 25514 14660 25570 14662
rect 21800 14170 21856 14172
rect 21880 14170 21936 14172
rect 21960 14170 22016 14172
rect 22040 14170 22096 14172
rect 21800 14118 21846 14170
rect 21846 14118 21856 14170
rect 21880 14118 21910 14170
rect 21910 14118 21922 14170
rect 21922 14118 21936 14170
rect 21960 14118 21974 14170
rect 21974 14118 21986 14170
rect 21986 14118 22016 14170
rect 22040 14118 22050 14170
rect 22050 14118 22096 14170
rect 21800 14116 21856 14118
rect 21880 14116 21936 14118
rect 21960 14116 22016 14118
rect 22040 14116 22096 14118
rect 18326 13626 18382 13628
rect 18406 13626 18462 13628
rect 18486 13626 18542 13628
rect 18566 13626 18622 13628
rect 18326 13574 18372 13626
rect 18372 13574 18382 13626
rect 18406 13574 18436 13626
rect 18436 13574 18448 13626
rect 18448 13574 18462 13626
rect 18486 13574 18500 13626
rect 18500 13574 18512 13626
rect 18512 13574 18542 13626
rect 18566 13574 18576 13626
rect 18576 13574 18622 13626
rect 18326 13572 18382 13574
rect 18406 13572 18462 13574
rect 18486 13572 18542 13574
rect 18566 13572 18622 13574
rect 25274 13626 25330 13628
rect 25354 13626 25410 13628
rect 25434 13626 25490 13628
rect 25514 13626 25570 13628
rect 25274 13574 25320 13626
rect 25320 13574 25330 13626
rect 25354 13574 25384 13626
rect 25384 13574 25396 13626
rect 25396 13574 25410 13626
rect 25434 13574 25448 13626
rect 25448 13574 25460 13626
rect 25460 13574 25490 13626
rect 25514 13574 25524 13626
rect 25524 13574 25570 13626
rect 25274 13572 25330 13574
rect 25354 13572 25410 13574
rect 25434 13572 25490 13574
rect 25514 13572 25570 13574
rect 21800 13082 21856 13084
rect 21880 13082 21936 13084
rect 21960 13082 22016 13084
rect 22040 13082 22096 13084
rect 21800 13030 21846 13082
rect 21846 13030 21856 13082
rect 21880 13030 21910 13082
rect 21910 13030 21922 13082
rect 21922 13030 21936 13082
rect 21960 13030 21974 13082
rect 21974 13030 21986 13082
rect 21986 13030 22016 13082
rect 22040 13030 22050 13082
rect 22050 13030 22096 13082
rect 21800 13028 21856 13030
rect 21880 13028 21936 13030
rect 21960 13028 22016 13030
rect 22040 13028 22096 13030
rect 18326 12538 18382 12540
rect 18406 12538 18462 12540
rect 18486 12538 18542 12540
rect 18566 12538 18622 12540
rect 18326 12486 18372 12538
rect 18372 12486 18382 12538
rect 18406 12486 18436 12538
rect 18436 12486 18448 12538
rect 18448 12486 18462 12538
rect 18486 12486 18500 12538
rect 18500 12486 18512 12538
rect 18512 12486 18542 12538
rect 18566 12486 18576 12538
rect 18576 12486 18622 12538
rect 18326 12484 18382 12486
rect 18406 12484 18462 12486
rect 18486 12484 18542 12486
rect 18566 12484 18622 12486
rect 25274 12538 25330 12540
rect 25354 12538 25410 12540
rect 25434 12538 25490 12540
rect 25514 12538 25570 12540
rect 25274 12486 25320 12538
rect 25320 12486 25330 12538
rect 25354 12486 25384 12538
rect 25384 12486 25396 12538
rect 25396 12486 25410 12538
rect 25434 12486 25448 12538
rect 25448 12486 25460 12538
rect 25460 12486 25490 12538
rect 25514 12486 25524 12538
rect 25524 12486 25570 12538
rect 25274 12484 25330 12486
rect 25354 12484 25410 12486
rect 25434 12484 25490 12486
rect 25514 12484 25570 12486
rect 21800 11994 21856 11996
rect 21880 11994 21936 11996
rect 21960 11994 22016 11996
rect 22040 11994 22096 11996
rect 21800 11942 21846 11994
rect 21846 11942 21856 11994
rect 21880 11942 21910 11994
rect 21910 11942 21922 11994
rect 21922 11942 21936 11994
rect 21960 11942 21974 11994
rect 21974 11942 21986 11994
rect 21986 11942 22016 11994
rect 22040 11942 22050 11994
rect 22050 11942 22096 11994
rect 21800 11940 21856 11942
rect 21880 11940 21936 11942
rect 21960 11940 22016 11942
rect 22040 11940 22096 11942
rect 18326 11450 18382 11452
rect 18406 11450 18462 11452
rect 18486 11450 18542 11452
rect 18566 11450 18622 11452
rect 18326 11398 18372 11450
rect 18372 11398 18382 11450
rect 18406 11398 18436 11450
rect 18436 11398 18448 11450
rect 18448 11398 18462 11450
rect 18486 11398 18500 11450
rect 18500 11398 18512 11450
rect 18512 11398 18542 11450
rect 18566 11398 18576 11450
rect 18576 11398 18622 11450
rect 18326 11396 18382 11398
rect 18406 11396 18462 11398
rect 18486 11396 18542 11398
rect 18566 11396 18622 11398
rect 25274 11450 25330 11452
rect 25354 11450 25410 11452
rect 25434 11450 25490 11452
rect 25514 11450 25570 11452
rect 25274 11398 25320 11450
rect 25320 11398 25330 11450
rect 25354 11398 25384 11450
rect 25384 11398 25396 11450
rect 25396 11398 25410 11450
rect 25434 11398 25448 11450
rect 25448 11398 25460 11450
rect 25460 11398 25490 11450
rect 25514 11398 25524 11450
rect 25524 11398 25570 11450
rect 25274 11396 25330 11398
rect 25354 11396 25410 11398
rect 25434 11396 25490 11398
rect 25514 11396 25570 11398
rect 21800 10906 21856 10908
rect 21880 10906 21936 10908
rect 21960 10906 22016 10908
rect 22040 10906 22096 10908
rect 21800 10854 21846 10906
rect 21846 10854 21856 10906
rect 21880 10854 21910 10906
rect 21910 10854 21922 10906
rect 21922 10854 21936 10906
rect 21960 10854 21974 10906
rect 21974 10854 21986 10906
rect 21986 10854 22016 10906
rect 22040 10854 22050 10906
rect 22050 10854 22096 10906
rect 21800 10852 21856 10854
rect 21880 10852 21936 10854
rect 21960 10852 22016 10854
rect 22040 10852 22096 10854
rect 18326 10362 18382 10364
rect 18406 10362 18462 10364
rect 18486 10362 18542 10364
rect 18566 10362 18622 10364
rect 18326 10310 18372 10362
rect 18372 10310 18382 10362
rect 18406 10310 18436 10362
rect 18436 10310 18448 10362
rect 18448 10310 18462 10362
rect 18486 10310 18500 10362
rect 18500 10310 18512 10362
rect 18512 10310 18542 10362
rect 18566 10310 18576 10362
rect 18576 10310 18622 10362
rect 18326 10308 18382 10310
rect 18406 10308 18462 10310
rect 18486 10308 18542 10310
rect 18566 10308 18622 10310
rect 25274 10362 25330 10364
rect 25354 10362 25410 10364
rect 25434 10362 25490 10364
rect 25514 10362 25570 10364
rect 25274 10310 25320 10362
rect 25320 10310 25330 10362
rect 25354 10310 25384 10362
rect 25384 10310 25396 10362
rect 25396 10310 25410 10362
rect 25434 10310 25448 10362
rect 25448 10310 25460 10362
rect 25460 10310 25490 10362
rect 25514 10310 25524 10362
rect 25524 10310 25570 10362
rect 25274 10308 25330 10310
rect 25354 10308 25410 10310
rect 25434 10308 25490 10310
rect 25514 10308 25570 10310
rect 21800 9818 21856 9820
rect 21880 9818 21936 9820
rect 21960 9818 22016 9820
rect 22040 9818 22096 9820
rect 21800 9766 21846 9818
rect 21846 9766 21856 9818
rect 21880 9766 21910 9818
rect 21910 9766 21922 9818
rect 21922 9766 21936 9818
rect 21960 9766 21974 9818
rect 21974 9766 21986 9818
rect 21986 9766 22016 9818
rect 22040 9766 22050 9818
rect 22050 9766 22096 9818
rect 21800 9764 21856 9766
rect 21880 9764 21936 9766
rect 21960 9764 22016 9766
rect 22040 9764 22096 9766
rect 18326 9274 18382 9276
rect 18406 9274 18462 9276
rect 18486 9274 18542 9276
rect 18566 9274 18622 9276
rect 18326 9222 18372 9274
rect 18372 9222 18382 9274
rect 18406 9222 18436 9274
rect 18436 9222 18448 9274
rect 18448 9222 18462 9274
rect 18486 9222 18500 9274
rect 18500 9222 18512 9274
rect 18512 9222 18542 9274
rect 18566 9222 18576 9274
rect 18576 9222 18622 9274
rect 18326 9220 18382 9222
rect 18406 9220 18462 9222
rect 18486 9220 18542 9222
rect 18566 9220 18622 9222
rect 18326 8186 18382 8188
rect 18406 8186 18462 8188
rect 18486 8186 18542 8188
rect 18566 8186 18622 8188
rect 18326 8134 18372 8186
rect 18372 8134 18382 8186
rect 18406 8134 18436 8186
rect 18436 8134 18448 8186
rect 18448 8134 18462 8186
rect 18486 8134 18500 8186
rect 18500 8134 18512 8186
rect 18512 8134 18542 8186
rect 18566 8134 18576 8186
rect 18576 8134 18622 8186
rect 18326 8132 18382 8134
rect 18406 8132 18462 8134
rect 18486 8132 18542 8134
rect 18566 8132 18622 8134
rect 18326 7098 18382 7100
rect 18406 7098 18462 7100
rect 18486 7098 18542 7100
rect 18566 7098 18622 7100
rect 18326 7046 18372 7098
rect 18372 7046 18382 7098
rect 18406 7046 18436 7098
rect 18436 7046 18448 7098
rect 18448 7046 18462 7098
rect 18486 7046 18500 7098
rect 18500 7046 18512 7098
rect 18512 7046 18542 7098
rect 18566 7046 18576 7098
rect 18576 7046 18622 7098
rect 18326 7044 18382 7046
rect 18406 7044 18462 7046
rect 18486 7044 18542 7046
rect 18566 7044 18622 7046
rect 25274 9274 25330 9276
rect 25354 9274 25410 9276
rect 25434 9274 25490 9276
rect 25514 9274 25570 9276
rect 25274 9222 25320 9274
rect 25320 9222 25330 9274
rect 25354 9222 25384 9274
rect 25384 9222 25396 9274
rect 25396 9222 25410 9274
rect 25434 9222 25448 9274
rect 25448 9222 25460 9274
rect 25460 9222 25490 9274
rect 25514 9222 25524 9274
rect 25524 9222 25570 9274
rect 25274 9220 25330 9222
rect 25354 9220 25410 9222
rect 25434 9220 25490 9222
rect 25514 9220 25570 9222
rect 21800 8730 21856 8732
rect 21880 8730 21936 8732
rect 21960 8730 22016 8732
rect 22040 8730 22096 8732
rect 21800 8678 21846 8730
rect 21846 8678 21856 8730
rect 21880 8678 21910 8730
rect 21910 8678 21922 8730
rect 21922 8678 21936 8730
rect 21960 8678 21974 8730
rect 21974 8678 21986 8730
rect 21986 8678 22016 8730
rect 22040 8678 22050 8730
rect 22050 8678 22096 8730
rect 21800 8676 21856 8678
rect 21880 8676 21936 8678
rect 21960 8676 22016 8678
rect 22040 8676 22096 8678
rect 25274 8186 25330 8188
rect 25354 8186 25410 8188
rect 25434 8186 25490 8188
rect 25514 8186 25570 8188
rect 25274 8134 25320 8186
rect 25320 8134 25330 8186
rect 25354 8134 25384 8186
rect 25384 8134 25396 8186
rect 25396 8134 25410 8186
rect 25434 8134 25448 8186
rect 25448 8134 25460 8186
rect 25460 8134 25490 8186
rect 25514 8134 25524 8186
rect 25524 8134 25570 8186
rect 25274 8132 25330 8134
rect 25354 8132 25410 8134
rect 25434 8132 25490 8134
rect 25514 8132 25570 8134
rect 21800 7642 21856 7644
rect 21880 7642 21936 7644
rect 21960 7642 22016 7644
rect 22040 7642 22096 7644
rect 21800 7590 21846 7642
rect 21846 7590 21856 7642
rect 21880 7590 21910 7642
rect 21910 7590 21922 7642
rect 21922 7590 21936 7642
rect 21960 7590 21974 7642
rect 21974 7590 21986 7642
rect 21986 7590 22016 7642
rect 22040 7590 22050 7642
rect 22050 7590 22096 7642
rect 21800 7588 21856 7590
rect 21880 7588 21936 7590
rect 21960 7588 22016 7590
rect 22040 7588 22096 7590
rect 14852 6554 14908 6556
rect 14932 6554 14988 6556
rect 15012 6554 15068 6556
rect 15092 6554 15148 6556
rect 14852 6502 14898 6554
rect 14898 6502 14908 6554
rect 14932 6502 14962 6554
rect 14962 6502 14974 6554
rect 14974 6502 14988 6554
rect 15012 6502 15026 6554
rect 15026 6502 15038 6554
rect 15038 6502 15068 6554
rect 15092 6502 15102 6554
rect 15102 6502 15148 6554
rect 14852 6500 14908 6502
rect 14932 6500 14988 6502
rect 15012 6500 15068 6502
rect 15092 6500 15148 6502
rect 18970 6704 19026 6760
rect 21800 6554 21856 6556
rect 21880 6554 21936 6556
rect 21960 6554 22016 6556
rect 22040 6554 22096 6556
rect 21800 6502 21846 6554
rect 21846 6502 21856 6554
rect 21880 6502 21910 6554
rect 21910 6502 21922 6554
rect 21922 6502 21936 6554
rect 21960 6502 21974 6554
rect 21974 6502 21986 6554
rect 21986 6502 22016 6554
rect 22040 6502 22050 6554
rect 22050 6502 22096 6554
rect 21800 6500 21856 6502
rect 21880 6500 21936 6502
rect 21960 6500 22016 6502
rect 22040 6500 22096 6502
rect 16578 6296 16634 6352
rect 14852 5466 14908 5468
rect 14932 5466 14988 5468
rect 15012 5466 15068 5468
rect 15092 5466 15148 5468
rect 14852 5414 14898 5466
rect 14898 5414 14908 5466
rect 14932 5414 14962 5466
rect 14962 5414 14974 5466
rect 14974 5414 14988 5466
rect 15012 5414 15026 5466
rect 15026 5414 15038 5466
rect 15038 5414 15068 5466
rect 15092 5414 15102 5466
rect 15102 5414 15148 5466
rect 14852 5412 14908 5414
rect 14932 5412 14988 5414
rect 15012 5412 15068 5414
rect 15092 5412 15148 5414
rect 18326 6010 18382 6012
rect 18406 6010 18462 6012
rect 18486 6010 18542 6012
rect 18566 6010 18622 6012
rect 18326 5958 18372 6010
rect 18372 5958 18382 6010
rect 18406 5958 18436 6010
rect 18436 5958 18448 6010
rect 18448 5958 18462 6010
rect 18486 5958 18500 6010
rect 18500 5958 18512 6010
rect 18512 5958 18542 6010
rect 18566 5958 18576 6010
rect 18576 5958 18622 6010
rect 18326 5956 18382 5958
rect 18406 5956 18462 5958
rect 18486 5956 18542 5958
rect 18566 5956 18622 5958
rect 21800 5466 21856 5468
rect 21880 5466 21936 5468
rect 21960 5466 22016 5468
rect 22040 5466 22096 5468
rect 21800 5414 21846 5466
rect 21846 5414 21856 5466
rect 21880 5414 21910 5466
rect 21910 5414 21922 5466
rect 21922 5414 21936 5466
rect 21960 5414 21974 5466
rect 21974 5414 21986 5466
rect 21986 5414 22016 5466
rect 22040 5414 22050 5466
rect 22050 5414 22096 5466
rect 21800 5412 21856 5414
rect 21880 5412 21936 5414
rect 21960 5412 22016 5414
rect 22040 5412 22096 5414
rect 18326 4922 18382 4924
rect 18406 4922 18462 4924
rect 18486 4922 18542 4924
rect 18566 4922 18622 4924
rect 18326 4870 18372 4922
rect 18372 4870 18382 4922
rect 18406 4870 18436 4922
rect 18436 4870 18448 4922
rect 18448 4870 18462 4922
rect 18486 4870 18500 4922
rect 18500 4870 18512 4922
rect 18512 4870 18542 4922
rect 18566 4870 18576 4922
rect 18576 4870 18622 4922
rect 18326 4868 18382 4870
rect 18406 4868 18462 4870
rect 18486 4868 18542 4870
rect 18566 4868 18622 4870
rect 14852 4378 14908 4380
rect 14932 4378 14988 4380
rect 15012 4378 15068 4380
rect 15092 4378 15148 4380
rect 14852 4326 14898 4378
rect 14898 4326 14908 4378
rect 14932 4326 14962 4378
rect 14962 4326 14974 4378
rect 14974 4326 14988 4378
rect 15012 4326 15026 4378
rect 15026 4326 15038 4378
rect 15038 4326 15068 4378
rect 15092 4326 15102 4378
rect 15102 4326 15148 4378
rect 14852 4324 14908 4326
rect 14932 4324 14988 4326
rect 15012 4324 15068 4326
rect 15092 4324 15148 4326
rect 14852 3290 14908 3292
rect 14932 3290 14988 3292
rect 15012 3290 15068 3292
rect 15092 3290 15148 3292
rect 14852 3238 14898 3290
rect 14898 3238 14908 3290
rect 14932 3238 14962 3290
rect 14962 3238 14974 3290
rect 14974 3238 14988 3290
rect 15012 3238 15026 3290
rect 15026 3238 15038 3290
rect 15038 3238 15068 3290
rect 15092 3238 15102 3290
rect 15102 3238 15148 3290
rect 14852 3236 14908 3238
rect 14932 3236 14988 3238
rect 15012 3236 15068 3238
rect 15092 3236 15148 3238
rect 11378 2746 11434 2748
rect 11458 2746 11514 2748
rect 11538 2746 11594 2748
rect 11618 2746 11674 2748
rect 11378 2694 11424 2746
rect 11424 2694 11434 2746
rect 11458 2694 11488 2746
rect 11488 2694 11500 2746
rect 11500 2694 11514 2746
rect 11538 2694 11552 2746
rect 11552 2694 11564 2746
rect 11564 2694 11594 2746
rect 11618 2694 11628 2746
rect 11628 2694 11674 2746
rect 11378 2692 11434 2694
rect 11458 2692 11514 2694
rect 11538 2692 11594 2694
rect 11618 2692 11674 2694
rect 21800 4378 21856 4380
rect 21880 4378 21936 4380
rect 21960 4378 22016 4380
rect 22040 4378 22096 4380
rect 21800 4326 21846 4378
rect 21846 4326 21856 4378
rect 21880 4326 21910 4378
rect 21910 4326 21922 4378
rect 21922 4326 21936 4378
rect 21960 4326 21974 4378
rect 21974 4326 21986 4378
rect 21986 4326 22016 4378
rect 22040 4326 22050 4378
rect 22050 4326 22096 4378
rect 21800 4324 21856 4326
rect 21880 4324 21936 4326
rect 21960 4324 22016 4326
rect 22040 4324 22096 4326
rect 18326 3834 18382 3836
rect 18406 3834 18462 3836
rect 18486 3834 18542 3836
rect 18566 3834 18622 3836
rect 18326 3782 18372 3834
rect 18372 3782 18382 3834
rect 18406 3782 18436 3834
rect 18436 3782 18448 3834
rect 18448 3782 18462 3834
rect 18486 3782 18500 3834
rect 18500 3782 18512 3834
rect 18512 3782 18542 3834
rect 18566 3782 18576 3834
rect 18576 3782 18622 3834
rect 18326 3780 18382 3782
rect 18406 3780 18462 3782
rect 18486 3780 18542 3782
rect 18566 3780 18622 3782
rect 21800 3290 21856 3292
rect 21880 3290 21936 3292
rect 21960 3290 22016 3292
rect 22040 3290 22096 3292
rect 21800 3238 21846 3290
rect 21846 3238 21856 3290
rect 21880 3238 21910 3290
rect 21910 3238 21922 3290
rect 21922 3238 21936 3290
rect 21960 3238 21974 3290
rect 21974 3238 21986 3290
rect 21986 3238 22016 3290
rect 22040 3238 22050 3290
rect 22050 3238 22096 3290
rect 21800 3236 21856 3238
rect 21880 3236 21936 3238
rect 21960 3236 22016 3238
rect 22040 3236 22096 3238
rect 18326 2746 18382 2748
rect 18406 2746 18462 2748
rect 18486 2746 18542 2748
rect 18566 2746 18622 2748
rect 18326 2694 18372 2746
rect 18372 2694 18382 2746
rect 18406 2694 18436 2746
rect 18436 2694 18448 2746
rect 18448 2694 18462 2746
rect 18486 2694 18500 2746
rect 18500 2694 18512 2746
rect 18512 2694 18542 2746
rect 18566 2694 18576 2746
rect 18576 2694 18622 2746
rect 18326 2692 18382 2694
rect 18406 2692 18462 2694
rect 18486 2692 18542 2694
rect 18566 2692 18622 2694
rect 25274 7098 25330 7100
rect 25354 7098 25410 7100
rect 25434 7098 25490 7100
rect 25514 7098 25570 7100
rect 25274 7046 25320 7098
rect 25320 7046 25330 7098
rect 25354 7046 25384 7098
rect 25384 7046 25396 7098
rect 25396 7046 25410 7098
rect 25434 7046 25448 7098
rect 25448 7046 25460 7098
rect 25460 7046 25490 7098
rect 25514 7046 25524 7098
rect 25524 7046 25570 7098
rect 25274 7044 25330 7046
rect 25354 7044 25410 7046
rect 25434 7044 25490 7046
rect 25514 7044 25570 7046
rect 25274 6010 25330 6012
rect 25354 6010 25410 6012
rect 25434 6010 25490 6012
rect 25514 6010 25570 6012
rect 25274 5958 25320 6010
rect 25320 5958 25330 6010
rect 25354 5958 25384 6010
rect 25384 5958 25396 6010
rect 25396 5958 25410 6010
rect 25434 5958 25448 6010
rect 25448 5958 25460 6010
rect 25460 5958 25490 6010
rect 25514 5958 25524 6010
rect 25524 5958 25570 6010
rect 25274 5956 25330 5958
rect 25354 5956 25410 5958
rect 25434 5956 25490 5958
rect 25514 5956 25570 5958
rect 25274 4922 25330 4924
rect 25354 4922 25410 4924
rect 25434 4922 25490 4924
rect 25514 4922 25570 4924
rect 25274 4870 25320 4922
rect 25320 4870 25330 4922
rect 25354 4870 25384 4922
rect 25384 4870 25396 4922
rect 25396 4870 25410 4922
rect 25434 4870 25448 4922
rect 25448 4870 25460 4922
rect 25460 4870 25490 4922
rect 25514 4870 25524 4922
rect 25524 4870 25570 4922
rect 25274 4868 25330 4870
rect 25354 4868 25410 4870
rect 25434 4868 25490 4870
rect 25514 4868 25570 4870
rect 25274 3834 25330 3836
rect 25354 3834 25410 3836
rect 25434 3834 25490 3836
rect 25514 3834 25570 3836
rect 25274 3782 25320 3834
rect 25320 3782 25330 3834
rect 25354 3782 25384 3834
rect 25384 3782 25396 3834
rect 25396 3782 25410 3834
rect 25434 3782 25448 3834
rect 25448 3782 25460 3834
rect 25460 3782 25490 3834
rect 25514 3782 25524 3834
rect 25524 3782 25570 3834
rect 25274 3780 25330 3782
rect 25354 3780 25410 3782
rect 25434 3780 25490 3782
rect 25514 3780 25570 3782
rect 25274 2746 25330 2748
rect 25354 2746 25410 2748
rect 25434 2746 25490 2748
rect 25514 2746 25570 2748
rect 25274 2694 25320 2746
rect 25320 2694 25330 2746
rect 25354 2694 25384 2746
rect 25384 2694 25396 2746
rect 25396 2694 25410 2746
rect 25434 2694 25448 2746
rect 25448 2694 25460 2746
rect 25460 2694 25490 2746
rect 25514 2694 25524 2746
rect 25524 2694 25570 2746
rect 25274 2692 25330 2694
rect 25354 2692 25410 2694
rect 25434 2692 25490 2694
rect 25514 2692 25570 2694
rect 7904 2202 7960 2204
rect 7984 2202 8040 2204
rect 8064 2202 8120 2204
rect 8144 2202 8200 2204
rect 7904 2150 7950 2202
rect 7950 2150 7960 2202
rect 7984 2150 8014 2202
rect 8014 2150 8026 2202
rect 8026 2150 8040 2202
rect 8064 2150 8078 2202
rect 8078 2150 8090 2202
rect 8090 2150 8120 2202
rect 8144 2150 8154 2202
rect 8154 2150 8200 2202
rect 7904 2148 7960 2150
rect 7984 2148 8040 2150
rect 8064 2148 8120 2150
rect 8144 2148 8200 2150
rect 14852 2202 14908 2204
rect 14932 2202 14988 2204
rect 15012 2202 15068 2204
rect 15092 2202 15148 2204
rect 14852 2150 14898 2202
rect 14898 2150 14908 2202
rect 14932 2150 14962 2202
rect 14962 2150 14974 2202
rect 14974 2150 14988 2202
rect 15012 2150 15026 2202
rect 15026 2150 15038 2202
rect 15038 2150 15068 2202
rect 15092 2150 15102 2202
rect 15102 2150 15148 2202
rect 14852 2148 14908 2150
rect 14932 2148 14988 2150
rect 15012 2148 15068 2150
rect 15092 2148 15148 2150
rect 21800 2202 21856 2204
rect 21880 2202 21936 2204
rect 21960 2202 22016 2204
rect 22040 2202 22096 2204
rect 21800 2150 21846 2202
rect 21846 2150 21856 2202
rect 21880 2150 21910 2202
rect 21910 2150 21922 2202
rect 21922 2150 21936 2202
rect 21960 2150 21974 2202
rect 21974 2150 21986 2202
rect 21986 2150 22016 2202
rect 22040 2150 22050 2202
rect 22050 2150 22096 2202
rect 21800 2148 21856 2150
rect 21880 2148 21936 2150
rect 21960 2148 22016 2150
rect 22040 2148 22096 2150
<< metal3 >>
rect 4420 27776 4736 27777
rect 4420 27712 4426 27776
rect 4490 27712 4506 27776
rect 4570 27712 4586 27776
rect 4650 27712 4666 27776
rect 4730 27712 4736 27776
rect 4420 27711 4736 27712
rect 11368 27776 11684 27777
rect 11368 27712 11374 27776
rect 11438 27712 11454 27776
rect 11518 27712 11534 27776
rect 11598 27712 11614 27776
rect 11678 27712 11684 27776
rect 11368 27711 11684 27712
rect 18316 27776 18632 27777
rect 18316 27712 18322 27776
rect 18386 27712 18402 27776
rect 18466 27712 18482 27776
rect 18546 27712 18562 27776
rect 18626 27712 18632 27776
rect 18316 27711 18632 27712
rect 25264 27776 25580 27777
rect 25264 27712 25270 27776
rect 25334 27712 25350 27776
rect 25414 27712 25430 27776
rect 25494 27712 25510 27776
rect 25574 27712 25580 27776
rect 25264 27711 25580 27712
rect 7894 27232 8210 27233
rect 7894 27168 7900 27232
rect 7964 27168 7980 27232
rect 8044 27168 8060 27232
rect 8124 27168 8140 27232
rect 8204 27168 8210 27232
rect 7894 27167 8210 27168
rect 14842 27232 15158 27233
rect 14842 27168 14848 27232
rect 14912 27168 14928 27232
rect 14992 27168 15008 27232
rect 15072 27168 15088 27232
rect 15152 27168 15158 27232
rect 14842 27167 15158 27168
rect 21790 27232 22106 27233
rect 21790 27168 21796 27232
rect 21860 27168 21876 27232
rect 21940 27168 21956 27232
rect 22020 27168 22036 27232
rect 22100 27168 22106 27232
rect 21790 27167 22106 27168
rect 4420 26688 4736 26689
rect 4420 26624 4426 26688
rect 4490 26624 4506 26688
rect 4570 26624 4586 26688
rect 4650 26624 4666 26688
rect 4730 26624 4736 26688
rect 4420 26623 4736 26624
rect 11368 26688 11684 26689
rect 11368 26624 11374 26688
rect 11438 26624 11454 26688
rect 11518 26624 11534 26688
rect 11598 26624 11614 26688
rect 11678 26624 11684 26688
rect 11368 26623 11684 26624
rect 18316 26688 18632 26689
rect 18316 26624 18322 26688
rect 18386 26624 18402 26688
rect 18466 26624 18482 26688
rect 18546 26624 18562 26688
rect 18626 26624 18632 26688
rect 18316 26623 18632 26624
rect 25264 26688 25580 26689
rect 25264 26624 25270 26688
rect 25334 26624 25350 26688
rect 25414 26624 25430 26688
rect 25494 26624 25510 26688
rect 25574 26624 25580 26688
rect 25264 26623 25580 26624
rect 7894 26144 8210 26145
rect 7894 26080 7900 26144
rect 7964 26080 7980 26144
rect 8044 26080 8060 26144
rect 8124 26080 8140 26144
rect 8204 26080 8210 26144
rect 7894 26079 8210 26080
rect 14842 26144 15158 26145
rect 14842 26080 14848 26144
rect 14912 26080 14928 26144
rect 14992 26080 15008 26144
rect 15072 26080 15088 26144
rect 15152 26080 15158 26144
rect 14842 26079 15158 26080
rect 21790 26144 22106 26145
rect 21790 26080 21796 26144
rect 21860 26080 21876 26144
rect 21940 26080 21956 26144
rect 22020 26080 22036 26144
rect 22100 26080 22106 26144
rect 21790 26079 22106 26080
rect 4420 25600 4736 25601
rect 4420 25536 4426 25600
rect 4490 25536 4506 25600
rect 4570 25536 4586 25600
rect 4650 25536 4666 25600
rect 4730 25536 4736 25600
rect 4420 25535 4736 25536
rect 11368 25600 11684 25601
rect 11368 25536 11374 25600
rect 11438 25536 11454 25600
rect 11518 25536 11534 25600
rect 11598 25536 11614 25600
rect 11678 25536 11684 25600
rect 11368 25535 11684 25536
rect 18316 25600 18632 25601
rect 18316 25536 18322 25600
rect 18386 25536 18402 25600
rect 18466 25536 18482 25600
rect 18546 25536 18562 25600
rect 18626 25536 18632 25600
rect 18316 25535 18632 25536
rect 25264 25600 25580 25601
rect 25264 25536 25270 25600
rect 25334 25536 25350 25600
rect 25414 25536 25430 25600
rect 25494 25536 25510 25600
rect 25574 25536 25580 25600
rect 25264 25535 25580 25536
rect 7894 25056 8210 25057
rect 7894 24992 7900 25056
rect 7964 24992 7980 25056
rect 8044 24992 8060 25056
rect 8124 24992 8140 25056
rect 8204 24992 8210 25056
rect 7894 24991 8210 24992
rect 14842 25056 15158 25057
rect 14842 24992 14848 25056
rect 14912 24992 14928 25056
rect 14992 24992 15008 25056
rect 15072 24992 15088 25056
rect 15152 24992 15158 25056
rect 14842 24991 15158 24992
rect 21790 25056 22106 25057
rect 21790 24992 21796 25056
rect 21860 24992 21876 25056
rect 21940 24992 21956 25056
rect 22020 24992 22036 25056
rect 22100 24992 22106 25056
rect 21790 24991 22106 24992
rect 0 24578 800 24608
rect 1485 24578 1551 24581
rect 0 24576 1551 24578
rect 0 24520 1490 24576
rect 1546 24520 1551 24576
rect 0 24518 1551 24520
rect 0 24488 800 24518
rect 1485 24515 1551 24518
rect 4420 24512 4736 24513
rect 4420 24448 4426 24512
rect 4490 24448 4506 24512
rect 4570 24448 4586 24512
rect 4650 24448 4666 24512
rect 4730 24448 4736 24512
rect 4420 24447 4736 24448
rect 11368 24512 11684 24513
rect 11368 24448 11374 24512
rect 11438 24448 11454 24512
rect 11518 24448 11534 24512
rect 11598 24448 11614 24512
rect 11678 24448 11684 24512
rect 11368 24447 11684 24448
rect 18316 24512 18632 24513
rect 18316 24448 18322 24512
rect 18386 24448 18402 24512
rect 18466 24448 18482 24512
rect 18546 24448 18562 24512
rect 18626 24448 18632 24512
rect 18316 24447 18632 24448
rect 25264 24512 25580 24513
rect 25264 24448 25270 24512
rect 25334 24448 25350 24512
rect 25414 24448 25430 24512
rect 25494 24448 25510 24512
rect 25574 24448 25580 24512
rect 25264 24447 25580 24448
rect 7894 23968 8210 23969
rect 7894 23904 7900 23968
rect 7964 23904 7980 23968
rect 8044 23904 8060 23968
rect 8124 23904 8140 23968
rect 8204 23904 8210 23968
rect 7894 23903 8210 23904
rect 14842 23968 15158 23969
rect 14842 23904 14848 23968
rect 14912 23904 14928 23968
rect 14992 23904 15008 23968
rect 15072 23904 15088 23968
rect 15152 23904 15158 23968
rect 14842 23903 15158 23904
rect 21790 23968 22106 23969
rect 21790 23904 21796 23968
rect 21860 23904 21876 23968
rect 21940 23904 21956 23968
rect 22020 23904 22036 23968
rect 22100 23904 22106 23968
rect 21790 23903 22106 23904
rect 4420 23424 4736 23425
rect 4420 23360 4426 23424
rect 4490 23360 4506 23424
rect 4570 23360 4586 23424
rect 4650 23360 4666 23424
rect 4730 23360 4736 23424
rect 4420 23359 4736 23360
rect 11368 23424 11684 23425
rect 11368 23360 11374 23424
rect 11438 23360 11454 23424
rect 11518 23360 11534 23424
rect 11598 23360 11614 23424
rect 11678 23360 11684 23424
rect 11368 23359 11684 23360
rect 18316 23424 18632 23425
rect 18316 23360 18322 23424
rect 18386 23360 18402 23424
rect 18466 23360 18482 23424
rect 18546 23360 18562 23424
rect 18626 23360 18632 23424
rect 18316 23359 18632 23360
rect 25264 23424 25580 23425
rect 25264 23360 25270 23424
rect 25334 23360 25350 23424
rect 25414 23360 25430 23424
rect 25494 23360 25510 23424
rect 25574 23360 25580 23424
rect 25264 23359 25580 23360
rect 7894 22880 8210 22881
rect 7894 22816 7900 22880
rect 7964 22816 7980 22880
rect 8044 22816 8060 22880
rect 8124 22816 8140 22880
rect 8204 22816 8210 22880
rect 7894 22815 8210 22816
rect 14842 22880 15158 22881
rect 14842 22816 14848 22880
rect 14912 22816 14928 22880
rect 14992 22816 15008 22880
rect 15072 22816 15088 22880
rect 15152 22816 15158 22880
rect 14842 22815 15158 22816
rect 21790 22880 22106 22881
rect 21790 22816 21796 22880
rect 21860 22816 21876 22880
rect 21940 22816 21956 22880
rect 22020 22816 22036 22880
rect 22100 22816 22106 22880
rect 21790 22815 22106 22816
rect 4420 22336 4736 22337
rect 4420 22272 4426 22336
rect 4490 22272 4506 22336
rect 4570 22272 4586 22336
rect 4650 22272 4666 22336
rect 4730 22272 4736 22336
rect 4420 22271 4736 22272
rect 11368 22336 11684 22337
rect 11368 22272 11374 22336
rect 11438 22272 11454 22336
rect 11518 22272 11534 22336
rect 11598 22272 11614 22336
rect 11678 22272 11684 22336
rect 11368 22271 11684 22272
rect 18316 22336 18632 22337
rect 18316 22272 18322 22336
rect 18386 22272 18402 22336
rect 18466 22272 18482 22336
rect 18546 22272 18562 22336
rect 18626 22272 18632 22336
rect 18316 22271 18632 22272
rect 25264 22336 25580 22337
rect 25264 22272 25270 22336
rect 25334 22272 25350 22336
rect 25414 22272 25430 22336
rect 25494 22272 25510 22336
rect 25574 22272 25580 22336
rect 25264 22271 25580 22272
rect 7894 21792 8210 21793
rect 7894 21728 7900 21792
rect 7964 21728 7980 21792
rect 8044 21728 8060 21792
rect 8124 21728 8140 21792
rect 8204 21728 8210 21792
rect 7894 21727 8210 21728
rect 14842 21792 15158 21793
rect 14842 21728 14848 21792
rect 14912 21728 14928 21792
rect 14992 21728 15008 21792
rect 15072 21728 15088 21792
rect 15152 21728 15158 21792
rect 14842 21727 15158 21728
rect 21790 21792 22106 21793
rect 21790 21728 21796 21792
rect 21860 21728 21876 21792
rect 21940 21728 21956 21792
rect 22020 21728 22036 21792
rect 22100 21728 22106 21792
rect 21790 21727 22106 21728
rect 4420 21248 4736 21249
rect 4420 21184 4426 21248
rect 4490 21184 4506 21248
rect 4570 21184 4586 21248
rect 4650 21184 4666 21248
rect 4730 21184 4736 21248
rect 4420 21183 4736 21184
rect 11368 21248 11684 21249
rect 11368 21184 11374 21248
rect 11438 21184 11454 21248
rect 11518 21184 11534 21248
rect 11598 21184 11614 21248
rect 11678 21184 11684 21248
rect 11368 21183 11684 21184
rect 18316 21248 18632 21249
rect 18316 21184 18322 21248
rect 18386 21184 18402 21248
rect 18466 21184 18482 21248
rect 18546 21184 18562 21248
rect 18626 21184 18632 21248
rect 18316 21183 18632 21184
rect 25264 21248 25580 21249
rect 25264 21184 25270 21248
rect 25334 21184 25350 21248
rect 25414 21184 25430 21248
rect 25494 21184 25510 21248
rect 25574 21184 25580 21248
rect 25264 21183 25580 21184
rect 7894 20704 8210 20705
rect 7894 20640 7900 20704
rect 7964 20640 7980 20704
rect 8044 20640 8060 20704
rect 8124 20640 8140 20704
rect 8204 20640 8210 20704
rect 7894 20639 8210 20640
rect 14842 20704 15158 20705
rect 14842 20640 14848 20704
rect 14912 20640 14928 20704
rect 14992 20640 15008 20704
rect 15072 20640 15088 20704
rect 15152 20640 15158 20704
rect 14842 20639 15158 20640
rect 21790 20704 22106 20705
rect 21790 20640 21796 20704
rect 21860 20640 21876 20704
rect 21940 20640 21956 20704
rect 22020 20640 22036 20704
rect 22100 20640 22106 20704
rect 21790 20639 22106 20640
rect 4420 20160 4736 20161
rect 4420 20096 4426 20160
rect 4490 20096 4506 20160
rect 4570 20096 4586 20160
rect 4650 20096 4666 20160
rect 4730 20096 4736 20160
rect 4420 20095 4736 20096
rect 11368 20160 11684 20161
rect 11368 20096 11374 20160
rect 11438 20096 11454 20160
rect 11518 20096 11534 20160
rect 11598 20096 11614 20160
rect 11678 20096 11684 20160
rect 11368 20095 11684 20096
rect 18316 20160 18632 20161
rect 18316 20096 18322 20160
rect 18386 20096 18402 20160
rect 18466 20096 18482 20160
rect 18546 20096 18562 20160
rect 18626 20096 18632 20160
rect 18316 20095 18632 20096
rect 25264 20160 25580 20161
rect 25264 20096 25270 20160
rect 25334 20096 25350 20160
rect 25414 20096 25430 20160
rect 25494 20096 25510 20160
rect 25574 20096 25580 20160
rect 25264 20095 25580 20096
rect 7894 19616 8210 19617
rect 7894 19552 7900 19616
rect 7964 19552 7980 19616
rect 8044 19552 8060 19616
rect 8124 19552 8140 19616
rect 8204 19552 8210 19616
rect 7894 19551 8210 19552
rect 14842 19616 15158 19617
rect 14842 19552 14848 19616
rect 14912 19552 14928 19616
rect 14992 19552 15008 19616
rect 15072 19552 15088 19616
rect 15152 19552 15158 19616
rect 14842 19551 15158 19552
rect 21790 19616 22106 19617
rect 21790 19552 21796 19616
rect 21860 19552 21876 19616
rect 21940 19552 21956 19616
rect 22020 19552 22036 19616
rect 22100 19552 22106 19616
rect 21790 19551 22106 19552
rect 4420 19072 4736 19073
rect 4420 19008 4426 19072
rect 4490 19008 4506 19072
rect 4570 19008 4586 19072
rect 4650 19008 4666 19072
rect 4730 19008 4736 19072
rect 4420 19007 4736 19008
rect 11368 19072 11684 19073
rect 11368 19008 11374 19072
rect 11438 19008 11454 19072
rect 11518 19008 11534 19072
rect 11598 19008 11614 19072
rect 11678 19008 11684 19072
rect 11368 19007 11684 19008
rect 18316 19072 18632 19073
rect 18316 19008 18322 19072
rect 18386 19008 18402 19072
rect 18466 19008 18482 19072
rect 18546 19008 18562 19072
rect 18626 19008 18632 19072
rect 18316 19007 18632 19008
rect 25264 19072 25580 19073
rect 25264 19008 25270 19072
rect 25334 19008 25350 19072
rect 25414 19008 25430 19072
rect 25494 19008 25510 19072
rect 25574 19008 25580 19072
rect 25264 19007 25580 19008
rect 7894 18528 8210 18529
rect 7894 18464 7900 18528
rect 7964 18464 7980 18528
rect 8044 18464 8060 18528
rect 8124 18464 8140 18528
rect 8204 18464 8210 18528
rect 7894 18463 8210 18464
rect 14842 18528 15158 18529
rect 14842 18464 14848 18528
rect 14912 18464 14928 18528
rect 14992 18464 15008 18528
rect 15072 18464 15088 18528
rect 15152 18464 15158 18528
rect 14842 18463 15158 18464
rect 21790 18528 22106 18529
rect 21790 18464 21796 18528
rect 21860 18464 21876 18528
rect 21940 18464 21956 18528
rect 22020 18464 22036 18528
rect 22100 18464 22106 18528
rect 21790 18463 22106 18464
rect 4420 17984 4736 17985
rect 4420 17920 4426 17984
rect 4490 17920 4506 17984
rect 4570 17920 4586 17984
rect 4650 17920 4666 17984
rect 4730 17920 4736 17984
rect 4420 17919 4736 17920
rect 11368 17984 11684 17985
rect 11368 17920 11374 17984
rect 11438 17920 11454 17984
rect 11518 17920 11534 17984
rect 11598 17920 11614 17984
rect 11678 17920 11684 17984
rect 11368 17919 11684 17920
rect 18316 17984 18632 17985
rect 18316 17920 18322 17984
rect 18386 17920 18402 17984
rect 18466 17920 18482 17984
rect 18546 17920 18562 17984
rect 18626 17920 18632 17984
rect 18316 17919 18632 17920
rect 25264 17984 25580 17985
rect 25264 17920 25270 17984
rect 25334 17920 25350 17984
rect 25414 17920 25430 17984
rect 25494 17920 25510 17984
rect 25574 17920 25580 17984
rect 25264 17919 25580 17920
rect 7894 17440 8210 17441
rect 7894 17376 7900 17440
rect 7964 17376 7980 17440
rect 8044 17376 8060 17440
rect 8124 17376 8140 17440
rect 8204 17376 8210 17440
rect 7894 17375 8210 17376
rect 14842 17440 15158 17441
rect 14842 17376 14848 17440
rect 14912 17376 14928 17440
rect 14992 17376 15008 17440
rect 15072 17376 15088 17440
rect 15152 17376 15158 17440
rect 14842 17375 15158 17376
rect 21790 17440 22106 17441
rect 21790 17376 21796 17440
rect 21860 17376 21876 17440
rect 21940 17376 21956 17440
rect 22020 17376 22036 17440
rect 22100 17376 22106 17440
rect 21790 17375 22106 17376
rect 28165 17098 28231 17101
rect 29200 17098 30000 17128
rect 28165 17096 30000 17098
rect 28165 17040 28170 17096
rect 28226 17040 30000 17096
rect 28165 17038 30000 17040
rect 28165 17035 28231 17038
rect 29200 17008 30000 17038
rect 4420 16896 4736 16897
rect 4420 16832 4426 16896
rect 4490 16832 4506 16896
rect 4570 16832 4586 16896
rect 4650 16832 4666 16896
rect 4730 16832 4736 16896
rect 4420 16831 4736 16832
rect 11368 16896 11684 16897
rect 11368 16832 11374 16896
rect 11438 16832 11454 16896
rect 11518 16832 11534 16896
rect 11598 16832 11614 16896
rect 11678 16832 11684 16896
rect 11368 16831 11684 16832
rect 18316 16896 18632 16897
rect 18316 16832 18322 16896
rect 18386 16832 18402 16896
rect 18466 16832 18482 16896
rect 18546 16832 18562 16896
rect 18626 16832 18632 16896
rect 18316 16831 18632 16832
rect 25264 16896 25580 16897
rect 25264 16832 25270 16896
rect 25334 16832 25350 16896
rect 25414 16832 25430 16896
rect 25494 16832 25510 16896
rect 25574 16832 25580 16896
rect 25264 16831 25580 16832
rect 7894 16352 8210 16353
rect 7894 16288 7900 16352
rect 7964 16288 7980 16352
rect 8044 16288 8060 16352
rect 8124 16288 8140 16352
rect 8204 16288 8210 16352
rect 7894 16287 8210 16288
rect 14842 16352 15158 16353
rect 14842 16288 14848 16352
rect 14912 16288 14928 16352
rect 14992 16288 15008 16352
rect 15072 16288 15088 16352
rect 15152 16288 15158 16352
rect 14842 16287 15158 16288
rect 21790 16352 22106 16353
rect 21790 16288 21796 16352
rect 21860 16288 21876 16352
rect 21940 16288 21956 16352
rect 22020 16288 22036 16352
rect 22100 16288 22106 16352
rect 21790 16287 22106 16288
rect 4420 15808 4736 15809
rect 4420 15744 4426 15808
rect 4490 15744 4506 15808
rect 4570 15744 4586 15808
rect 4650 15744 4666 15808
rect 4730 15744 4736 15808
rect 4420 15743 4736 15744
rect 11368 15808 11684 15809
rect 11368 15744 11374 15808
rect 11438 15744 11454 15808
rect 11518 15744 11534 15808
rect 11598 15744 11614 15808
rect 11678 15744 11684 15808
rect 11368 15743 11684 15744
rect 18316 15808 18632 15809
rect 18316 15744 18322 15808
rect 18386 15744 18402 15808
rect 18466 15744 18482 15808
rect 18546 15744 18562 15808
rect 18626 15744 18632 15808
rect 18316 15743 18632 15744
rect 25264 15808 25580 15809
rect 25264 15744 25270 15808
rect 25334 15744 25350 15808
rect 25414 15744 25430 15808
rect 25494 15744 25510 15808
rect 25574 15744 25580 15808
rect 25264 15743 25580 15744
rect 7894 15264 8210 15265
rect 7894 15200 7900 15264
rect 7964 15200 7980 15264
rect 8044 15200 8060 15264
rect 8124 15200 8140 15264
rect 8204 15200 8210 15264
rect 7894 15199 8210 15200
rect 14842 15264 15158 15265
rect 14842 15200 14848 15264
rect 14912 15200 14928 15264
rect 14992 15200 15008 15264
rect 15072 15200 15088 15264
rect 15152 15200 15158 15264
rect 14842 15199 15158 15200
rect 21790 15264 22106 15265
rect 21790 15200 21796 15264
rect 21860 15200 21876 15264
rect 21940 15200 21956 15264
rect 22020 15200 22036 15264
rect 22100 15200 22106 15264
rect 21790 15199 22106 15200
rect 4420 14720 4736 14721
rect 4420 14656 4426 14720
rect 4490 14656 4506 14720
rect 4570 14656 4586 14720
rect 4650 14656 4666 14720
rect 4730 14656 4736 14720
rect 4420 14655 4736 14656
rect 11368 14720 11684 14721
rect 11368 14656 11374 14720
rect 11438 14656 11454 14720
rect 11518 14656 11534 14720
rect 11598 14656 11614 14720
rect 11678 14656 11684 14720
rect 11368 14655 11684 14656
rect 18316 14720 18632 14721
rect 18316 14656 18322 14720
rect 18386 14656 18402 14720
rect 18466 14656 18482 14720
rect 18546 14656 18562 14720
rect 18626 14656 18632 14720
rect 18316 14655 18632 14656
rect 25264 14720 25580 14721
rect 25264 14656 25270 14720
rect 25334 14656 25350 14720
rect 25414 14656 25430 14720
rect 25494 14656 25510 14720
rect 25574 14656 25580 14720
rect 25264 14655 25580 14656
rect 7894 14176 8210 14177
rect 7894 14112 7900 14176
rect 7964 14112 7980 14176
rect 8044 14112 8060 14176
rect 8124 14112 8140 14176
rect 8204 14112 8210 14176
rect 7894 14111 8210 14112
rect 14842 14176 15158 14177
rect 14842 14112 14848 14176
rect 14912 14112 14928 14176
rect 14992 14112 15008 14176
rect 15072 14112 15088 14176
rect 15152 14112 15158 14176
rect 14842 14111 15158 14112
rect 21790 14176 22106 14177
rect 21790 14112 21796 14176
rect 21860 14112 21876 14176
rect 21940 14112 21956 14176
rect 22020 14112 22036 14176
rect 22100 14112 22106 14176
rect 21790 14111 22106 14112
rect 4420 13632 4736 13633
rect 4420 13568 4426 13632
rect 4490 13568 4506 13632
rect 4570 13568 4586 13632
rect 4650 13568 4666 13632
rect 4730 13568 4736 13632
rect 4420 13567 4736 13568
rect 11368 13632 11684 13633
rect 11368 13568 11374 13632
rect 11438 13568 11454 13632
rect 11518 13568 11534 13632
rect 11598 13568 11614 13632
rect 11678 13568 11684 13632
rect 11368 13567 11684 13568
rect 18316 13632 18632 13633
rect 18316 13568 18322 13632
rect 18386 13568 18402 13632
rect 18466 13568 18482 13632
rect 18546 13568 18562 13632
rect 18626 13568 18632 13632
rect 18316 13567 18632 13568
rect 25264 13632 25580 13633
rect 25264 13568 25270 13632
rect 25334 13568 25350 13632
rect 25414 13568 25430 13632
rect 25494 13568 25510 13632
rect 25574 13568 25580 13632
rect 25264 13567 25580 13568
rect 4245 13290 4311 13293
rect 11145 13290 11211 13293
rect 4245 13288 11211 13290
rect 4245 13232 4250 13288
rect 4306 13232 11150 13288
rect 11206 13232 11211 13288
rect 4245 13230 11211 13232
rect 4245 13227 4311 13230
rect 11145 13227 11211 13230
rect 7894 13088 8210 13089
rect 7894 13024 7900 13088
rect 7964 13024 7980 13088
rect 8044 13024 8060 13088
rect 8124 13024 8140 13088
rect 8204 13024 8210 13088
rect 7894 13023 8210 13024
rect 14842 13088 15158 13089
rect 14842 13024 14848 13088
rect 14912 13024 14928 13088
rect 14992 13024 15008 13088
rect 15072 13024 15088 13088
rect 15152 13024 15158 13088
rect 14842 13023 15158 13024
rect 21790 13088 22106 13089
rect 21790 13024 21796 13088
rect 21860 13024 21876 13088
rect 21940 13024 21956 13088
rect 22020 13024 22036 13088
rect 22100 13024 22106 13088
rect 21790 13023 22106 13024
rect 4420 12544 4736 12545
rect 4420 12480 4426 12544
rect 4490 12480 4506 12544
rect 4570 12480 4586 12544
rect 4650 12480 4666 12544
rect 4730 12480 4736 12544
rect 4420 12479 4736 12480
rect 11368 12544 11684 12545
rect 11368 12480 11374 12544
rect 11438 12480 11454 12544
rect 11518 12480 11534 12544
rect 11598 12480 11614 12544
rect 11678 12480 11684 12544
rect 11368 12479 11684 12480
rect 18316 12544 18632 12545
rect 18316 12480 18322 12544
rect 18386 12480 18402 12544
rect 18466 12480 18482 12544
rect 18546 12480 18562 12544
rect 18626 12480 18632 12544
rect 18316 12479 18632 12480
rect 25264 12544 25580 12545
rect 25264 12480 25270 12544
rect 25334 12480 25350 12544
rect 25414 12480 25430 12544
rect 25494 12480 25510 12544
rect 25574 12480 25580 12544
rect 25264 12479 25580 12480
rect 7894 12000 8210 12001
rect 7894 11936 7900 12000
rect 7964 11936 7980 12000
rect 8044 11936 8060 12000
rect 8124 11936 8140 12000
rect 8204 11936 8210 12000
rect 7894 11935 8210 11936
rect 14842 12000 15158 12001
rect 14842 11936 14848 12000
rect 14912 11936 14928 12000
rect 14992 11936 15008 12000
rect 15072 11936 15088 12000
rect 15152 11936 15158 12000
rect 14842 11935 15158 11936
rect 21790 12000 22106 12001
rect 21790 11936 21796 12000
rect 21860 11936 21876 12000
rect 21940 11936 21956 12000
rect 22020 11936 22036 12000
rect 22100 11936 22106 12000
rect 21790 11935 22106 11936
rect 4420 11456 4736 11457
rect 4420 11392 4426 11456
rect 4490 11392 4506 11456
rect 4570 11392 4586 11456
rect 4650 11392 4666 11456
rect 4730 11392 4736 11456
rect 4420 11391 4736 11392
rect 11368 11456 11684 11457
rect 11368 11392 11374 11456
rect 11438 11392 11454 11456
rect 11518 11392 11534 11456
rect 11598 11392 11614 11456
rect 11678 11392 11684 11456
rect 11368 11391 11684 11392
rect 18316 11456 18632 11457
rect 18316 11392 18322 11456
rect 18386 11392 18402 11456
rect 18466 11392 18482 11456
rect 18546 11392 18562 11456
rect 18626 11392 18632 11456
rect 18316 11391 18632 11392
rect 25264 11456 25580 11457
rect 25264 11392 25270 11456
rect 25334 11392 25350 11456
rect 25414 11392 25430 11456
rect 25494 11392 25510 11456
rect 25574 11392 25580 11456
rect 25264 11391 25580 11392
rect 7894 10912 8210 10913
rect 7894 10848 7900 10912
rect 7964 10848 7980 10912
rect 8044 10848 8060 10912
rect 8124 10848 8140 10912
rect 8204 10848 8210 10912
rect 7894 10847 8210 10848
rect 14842 10912 15158 10913
rect 14842 10848 14848 10912
rect 14912 10848 14928 10912
rect 14992 10848 15008 10912
rect 15072 10848 15088 10912
rect 15152 10848 15158 10912
rect 14842 10847 15158 10848
rect 21790 10912 22106 10913
rect 21790 10848 21796 10912
rect 21860 10848 21876 10912
rect 21940 10848 21956 10912
rect 22020 10848 22036 10912
rect 22100 10848 22106 10912
rect 21790 10847 22106 10848
rect 4420 10368 4736 10369
rect 4420 10304 4426 10368
rect 4490 10304 4506 10368
rect 4570 10304 4586 10368
rect 4650 10304 4666 10368
rect 4730 10304 4736 10368
rect 4420 10303 4736 10304
rect 11368 10368 11684 10369
rect 11368 10304 11374 10368
rect 11438 10304 11454 10368
rect 11518 10304 11534 10368
rect 11598 10304 11614 10368
rect 11678 10304 11684 10368
rect 11368 10303 11684 10304
rect 18316 10368 18632 10369
rect 18316 10304 18322 10368
rect 18386 10304 18402 10368
rect 18466 10304 18482 10368
rect 18546 10304 18562 10368
rect 18626 10304 18632 10368
rect 18316 10303 18632 10304
rect 25264 10368 25580 10369
rect 25264 10304 25270 10368
rect 25334 10304 25350 10368
rect 25414 10304 25430 10368
rect 25494 10304 25510 10368
rect 25574 10304 25580 10368
rect 25264 10303 25580 10304
rect 7894 9824 8210 9825
rect 7894 9760 7900 9824
rect 7964 9760 7980 9824
rect 8044 9760 8060 9824
rect 8124 9760 8140 9824
rect 8204 9760 8210 9824
rect 7894 9759 8210 9760
rect 14842 9824 15158 9825
rect 14842 9760 14848 9824
rect 14912 9760 14928 9824
rect 14992 9760 15008 9824
rect 15072 9760 15088 9824
rect 15152 9760 15158 9824
rect 14842 9759 15158 9760
rect 21790 9824 22106 9825
rect 21790 9760 21796 9824
rect 21860 9760 21876 9824
rect 21940 9760 21956 9824
rect 22020 9760 22036 9824
rect 22100 9760 22106 9824
rect 21790 9759 22106 9760
rect 4420 9280 4736 9281
rect 4420 9216 4426 9280
rect 4490 9216 4506 9280
rect 4570 9216 4586 9280
rect 4650 9216 4666 9280
rect 4730 9216 4736 9280
rect 4420 9215 4736 9216
rect 11368 9280 11684 9281
rect 11368 9216 11374 9280
rect 11438 9216 11454 9280
rect 11518 9216 11534 9280
rect 11598 9216 11614 9280
rect 11678 9216 11684 9280
rect 11368 9215 11684 9216
rect 18316 9280 18632 9281
rect 18316 9216 18322 9280
rect 18386 9216 18402 9280
rect 18466 9216 18482 9280
rect 18546 9216 18562 9280
rect 18626 9216 18632 9280
rect 18316 9215 18632 9216
rect 25264 9280 25580 9281
rect 25264 9216 25270 9280
rect 25334 9216 25350 9280
rect 25414 9216 25430 9280
rect 25494 9216 25510 9280
rect 25574 9216 25580 9280
rect 25264 9215 25580 9216
rect 7894 8736 8210 8737
rect 7894 8672 7900 8736
rect 7964 8672 7980 8736
rect 8044 8672 8060 8736
rect 8124 8672 8140 8736
rect 8204 8672 8210 8736
rect 7894 8671 8210 8672
rect 14842 8736 15158 8737
rect 14842 8672 14848 8736
rect 14912 8672 14928 8736
rect 14992 8672 15008 8736
rect 15072 8672 15088 8736
rect 15152 8672 15158 8736
rect 14842 8671 15158 8672
rect 21790 8736 22106 8737
rect 21790 8672 21796 8736
rect 21860 8672 21876 8736
rect 21940 8672 21956 8736
rect 22020 8672 22036 8736
rect 22100 8672 22106 8736
rect 21790 8671 22106 8672
rect 4420 8192 4736 8193
rect 4420 8128 4426 8192
rect 4490 8128 4506 8192
rect 4570 8128 4586 8192
rect 4650 8128 4666 8192
rect 4730 8128 4736 8192
rect 4420 8127 4736 8128
rect 11368 8192 11684 8193
rect 11368 8128 11374 8192
rect 11438 8128 11454 8192
rect 11518 8128 11534 8192
rect 11598 8128 11614 8192
rect 11678 8128 11684 8192
rect 11368 8127 11684 8128
rect 18316 8192 18632 8193
rect 18316 8128 18322 8192
rect 18386 8128 18402 8192
rect 18466 8128 18482 8192
rect 18546 8128 18562 8192
rect 18626 8128 18632 8192
rect 18316 8127 18632 8128
rect 25264 8192 25580 8193
rect 25264 8128 25270 8192
rect 25334 8128 25350 8192
rect 25414 8128 25430 8192
rect 25494 8128 25510 8192
rect 25574 8128 25580 8192
rect 25264 8127 25580 8128
rect 7894 7648 8210 7649
rect 7894 7584 7900 7648
rect 7964 7584 7980 7648
rect 8044 7584 8060 7648
rect 8124 7584 8140 7648
rect 8204 7584 8210 7648
rect 7894 7583 8210 7584
rect 14842 7648 15158 7649
rect 14842 7584 14848 7648
rect 14912 7584 14928 7648
rect 14992 7584 15008 7648
rect 15072 7584 15088 7648
rect 15152 7584 15158 7648
rect 14842 7583 15158 7584
rect 21790 7648 22106 7649
rect 21790 7584 21796 7648
rect 21860 7584 21876 7648
rect 21940 7584 21956 7648
rect 22020 7584 22036 7648
rect 22100 7584 22106 7648
rect 21790 7583 22106 7584
rect 4420 7104 4736 7105
rect 4420 7040 4426 7104
rect 4490 7040 4506 7104
rect 4570 7040 4586 7104
rect 4650 7040 4666 7104
rect 4730 7040 4736 7104
rect 4420 7039 4736 7040
rect 11368 7104 11684 7105
rect 11368 7040 11374 7104
rect 11438 7040 11454 7104
rect 11518 7040 11534 7104
rect 11598 7040 11614 7104
rect 11678 7040 11684 7104
rect 11368 7039 11684 7040
rect 18316 7104 18632 7105
rect 18316 7040 18322 7104
rect 18386 7040 18402 7104
rect 18466 7040 18482 7104
rect 18546 7040 18562 7104
rect 18626 7040 18632 7104
rect 18316 7039 18632 7040
rect 25264 7104 25580 7105
rect 25264 7040 25270 7104
rect 25334 7040 25350 7104
rect 25414 7040 25430 7104
rect 25494 7040 25510 7104
rect 25574 7040 25580 7104
rect 25264 7039 25580 7040
rect 5901 6898 5967 6901
rect 14089 6898 14155 6901
rect 5901 6896 14155 6898
rect 5901 6840 5906 6896
rect 5962 6840 14094 6896
rect 14150 6840 14155 6896
rect 5901 6838 14155 6840
rect 5901 6835 5967 6838
rect 14089 6835 14155 6838
rect 7741 6762 7807 6765
rect 18965 6762 19031 6765
rect 7741 6760 19031 6762
rect 7741 6704 7746 6760
rect 7802 6704 18970 6760
rect 19026 6704 19031 6760
rect 7741 6702 19031 6704
rect 7741 6699 7807 6702
rect 18965 6699 19031 6702
rect 7894 6560 8210 6561
rect 7894 6496 7900 6560
rect 7964 6496 7980 6560
rect 8044 6496 8060 6560
rect 8124 6496 8140 6560
rect 8204 6496 8210 6560
rect 7894 6495 8210 6496
rect 14842 6560 15158 6561
rect 14842 6496 14848 6560
rect 14912 6496 14928 6560
rect 14992 6496 15008 6560
rect 15072 6496 15088 6560
rect 15152 6496 15158 6560
rect 14842 6495 15158 6496
rect 21790 6560 22106 6561
rect 21790 6496 21796 6560
rect 21860 6496 21876 6560
rect 21940 6496 21956 6560
rect 22020 6496 22036 6560
rect 22100 6496 22106 6560
rect 21790 6495 22106 6496
rect 5349 6354 5415 6357
rect 16573 6354 16639 6357
rect 5349 6352 16639 6354
rect 5349 6296 5354 6352
rect 5410 6296 16578 6352
rect 16634 6296 16639 6352
rect 5349 6294 16639 6296
rect 5349 6291 5415 6294
rect 16573 6291 16639 6294
rect 4420 6016 4736 6017
rect 4420 5952 4426 6016
rect 4490 5952 4506 6016
rect 4570 5952 4586 6016
rect 4650 5952 4666 6016
rect 4730 5952 4736 6016
rect 4420 5951 4736 5952
rect 11368 6016 11684 6017
rect 11368 5952 11374 6016
rect 11438 5952 11454 6016
rect 11518 5952 11534 6016
rect 11598 5952 11614 6016
rect 11678 5952 11684 6016
rect 11368 5951 11684 5952
rect 18316 6016 18632 6017
rect 18316 5952 18322 6016
rect 18386 5952 18402 6016
rect 18466 5952 18482 6016
rect 18546 5952 18562 6016
rect 18626 5952 18632 6016
rect 18316 5951 18632 5952
rect 25264 6016 25580 6017
rect 25264 5952 25270 6016
rect 25334 5952 25350 6016
rect 25414 5952 25430 6016
rect 25494 5952 25510 6016
rect 25574 5952 25580 6016
rect 25264 5951 25580 5952
rect 7894 5472 8210 5473
rect 7894 5408 7900 5472
rect 7964 5408 7980 5472
rect 8044 5408 8060 5472
rect 8124 5408 8140 5472
rect 8204 5408 8210 5472
rect 7894 5407 8210 5408
rect 14842 5472 15158 5473
rect 14842 5408 14848 5472
rect 14912 5408 14928 5472
rect 14992 5408 15008 5472
rect 15072 5408 15088 5472
rect 15152 5408 15158 5472
rect 14842 5407 15158 5408
rect 21790 5472 22106 5473
rect 21790 5408 21796 5472
rect 21860 5408 21876 5472
rect 21940 5408 21956 5472
rect 22020 5408 22036 5472
rect 22100 5408 22106 5472
rect 21790 5407 22106 5408
rect 4420 4928 4736 4929
rect 4420 4864 4426 4928
rect 4490 4864 4506 4928
rect 4570 4864 4586 4928
rect 4650 4864 4666 4928
rect 4730 4864 4736 4928
rect 4420 4863 4736 4864
rect 11368 4928 11684 4929
rect 11368 4864 11374 4928
rect 11438 4864 11454 4928
rect 11518 4864 11534 4928
rect 11598 4864 11614 4928
rect 11678 4864 11684 4928
rect 11368 4863 11684 4864
rect 18316 4928 18632 4929
rect 18316 4864 18322 4928
rect 18386 4864 18402 4928
rect 18466 4864 18482 4928
rect 18546 4864 18562 4928
rect 18626 4864 18632 4928
rect 18316 4863 18632 4864
rect 25264 4928 25580 4929
rect 25264 4864 25270 4928
rect 25334 4864 25350 4928
rect 25414 4864 25430 4928
rect 25494 4864 25510 4928
rect 25574 4864 25580 4928
rect 25264 4863 25580 4864
rect 7894 4384 8210 4385
rect 7894 4320 7900 4384
rect 7964 4320 7980 4384
rect 8044 4320 8060 4384
rect 8124 4320 8140 4384
rect 8204 4320 8210 4384
rect 7894 4319 8210 4320
rect 14842 4384 15158 4385
rect 14842 4320 14848 4384
rect 14912 4320 14928 4384
rect 14992 4320 15008 4384
rect 15072 4320 15088 4384
rect 15152 4320 15158 4384
rect 14842 4319 15158 4320
rect 21790 4384 22106 4385
rect 21790 4320 21796 4384
rect 21860 4320 21876 4384
rect 21940 4320 21956 4384
rect 22020 4320 22036 4384
rect 22100 4320 22106 4384
rect 21790 4319 22106 4320
rect 4420 3840 4736 3841
rect 4420 3776 4426 3840
rect 4490 3776 4506 3840
rect 4570 3776 4586 3840
rect 4650 3776 4666 3840
rect 4730 3776 4736 3840
rect 4420 3775 4736 3776
rect 11368 3840 11684 3841
rect 11368 3776 11374 3840
rect 11438 3776 11454 3840
rect 11518 3776 11534 3840
rect 11598 3776 11614 3840
rect 11678 3776 11684 3840
rect 11368 3775 11684 3776
rect 18316 3840 18632 3841
rect 18316 3776 18322 3840
rect 18386 3776 18402 3840
rect 18466 3776 18482 3840
rect 18546 3776 18562 3840
rect 18626 3776 18632 3840
rect 18316 3775 18632 3776
rect 25264 3840 25580 3841
rect 25264 3776 25270 3840
rect 25334 3776 25350 3840
rect 25414 3776 25430 3840
rect 25494 3776 25510 3840
rect 25574 3776 25580 3840
rect 25264 3775 25580 3776
rect 7894 3296 8210 3297
rect 7894 3232 7900 3296
rect 7964 3232 7980 3296
rect 8044 3232 8060 3296
rect 8124 3232 8140 3296
rect 8204 3232 8210 3296
rect 7894 3231 8210 3232
rect 14842 3296 15158 3297
rect 14842 3232 14848 3296
rect 14912 3232 14928 3296
rect 14992 3232 15008 3296
rect 15072 3232 15088 3296
rect 15152 3232 15158 3296
rect 14842 3231 15158 3232
rect 21790 3296 22106 3297
rect 21790 3232 21796 3296
rect 21860 3232 21876 3296
rect 21940 3232 21956 3296
rect 22020 3232 22036 3296
rect 22100 3232 22106 3296
rect 21790 3231 22106 3232
rect 4420 2752 4736 2753
rect 4420 2688 4426 2752
rect 4490 2688 4506 2752
rect 4570 2688 4586 2752
rect 4650 2688 4666 2752
rect 4730 2688 4736 2752
rect 4420 2687 4736 2688
rect 11368 2752 11684 2753
rect 11368 2688 11374 2752
rect 11438 2688 11454 2752
rect 11518 2688 11534 2752
rect 11598 2688 11614 2752
rect 11678 2688 11684 2752
rect 11368 2687 11684 2688
rect 18316 2752 18632 2753
rect 18316 2688 18322 2752
rect 18386 2688 18402 2752
rect 18466 2688 18482 2752
rect 18546 2688 18562 2752
rect 18626 2688 18632 2752
rect 18316 2687 18632 2688
rect 25264 2752 25580 2753
rect 25264 2688 25270 2752
rect 25334 2688 25350 2752
rect 25414 2688 25430 2752
rect 25494 2688 25510 2752
rect 25574 2688 25580 2752
rect 25264 2687 25580 2688
rect 7894 2208 8210 2209
rect 7894 2144 7900 2208
rect 7964 2144 7980 2208
rect 8044 2144 8060 2208
rect 8124 2144 8140 2208
rect 8204 2144 8210 2208
rect 7894 2143 8210 2144
rect 14842 2208 15158 2209
rect 14842 2144 14848 2208
rect 14912 2144 14928 2208
rect 14992 2144 15008 2208
rect 15072 2144 15088 2208
rect 15152 2144 15158 2208
rect 14842 2143 15158 2144
rect 21790 2208 22106 2209
rect 21790 2144 21796 2208
rect 21860 2144 21876 2208
rect 21940 2144 21956 2208
rect 22020 2144 22036 2208
rect 22100 2144 22106 2208
rect 21790 2143 22106 2144
<< via3 >>
rect 4426 27772 4490 27776
rect 4426 27716 4430 27772
rect 4430 27716 4486 27772
rect 4486 27716 4490 27772
rect 4426 27712 4490 27716
rect 4506 27772 4570 27776
rect 4506 27716 4510 27772
rect 4510 27716 4566 27772
rect 4566 27716 4570 27772
rect 4506 27712 4570 27716
rect 4586 27772 4650 27776
rect 4586 27716 4590 27772
rect 4590 27716 4646 27772
rect 4646 27716 4650 27772
rect 4586 27712 4650 27716
rect 4666 27772 4730 27776
rect 4666 27716 4670 27772
rect 4670 27716 4726 27772
rect 4726 27716 4730 27772
rect 4666 27712 4730 27716
rect 11374 27772 11438 27776
rect 11374 27716 11378 27772
rect 11378 27716 11434 27772
rect 11434 27716 11438 27772
rect 11374 27712 11438 27716
rect 11454 27772 11518 27776
rect 11454 27716 11458 27772
rect 11458 27716 11514 27772
rect 11514 27716 11518 27772
rect 11454 27712 11518 27716
rect 11534 27772 11598 27776
rect 11534 27716 11538 27772
rect 11538 27716 11594 27772
rect 11594 27716 11598 27772
rect 11534 27712 11598 27716
rect 11614 27772 11678 27776
rect 11614 27716 11618 27772
rect 11618 27716 11674 27772
rect 11674 27716 11678 27772
rect 11614 27712 11678 27716
rect 18322 27772 18386 27776
rect 18322 27716 18326 27772
rect 18326 27716 18382 27772
rect 18382 27716 18386 27772
rect 18322 27712 18386 27716
rect 18402 27772 18466 27776
rect 18402 27716 18406 27772
rect 18406 27716 18462 27772
rect 18462 27716 18466 27772
rect 18402 27712 18466 27716
rect 18482 27772 18546 27776
rect 18482 27716 18486 27772
rect 18486 27716 18542 27772
rect 18542 27716 18546 27772
rect 18482 27712 18546 27716
rect 18562 27772 18626 27776
rect 18562 27716 18566 27772
rect 18566 27716 18622 27772
rect 18622 27716 18626 27772
rect 18562 27712 18626 27716
rect 25270 27772 25334 27776
rect 25270 27716 25274 27772
rect 25274 27716 25330 27772
rect 25330 27716 25334 27772
rect 25270 27712 25334 27716
rect 25350 27772 25414 27776
rect 25350 27716 25354 27772
rect 25354 27716 25410 27772
rect 25410 27716 25414 27772
rect 25350 27712 25414 27716
rect 25430 27772 25494 27776
rect 25430 27716 25434 27772
rect 25434 27716 25490 27772
rect 25490 27716 25494 27772
rect 25430 27712 25494 27716
rect 25510 27772 25574 27776
rect 25510 27716 25514 27772
rect 25514 27716 25570 27772
rect 25570 27716 25574 27772
rect 25510 27712 25574 27716
rect 7900 27228 7964 27232
rect 7900 27172 7904 27228
rect 7904 27172 7960 27228
rect 7960 27172 7964 27228
rect 7900 27168 7964 27172
rect 7980 27228 8044 27232
rect 7980 27172 7984 27228
rect 7984 27172 8040 27228
rect 8040 27172 8044 27228
rect 7980 27168 8044 27172
rect 8060 27228 8124 27232
rect 8060 27172 8064 27228
rect 8064 27172 8120 27228
rect 8120 27172 8124 27228
rect 8060 27168 8124 27172
rect 8140 27228 8204 27232
rect 8140 27172 8144 27228
rect 8144 27172 8200 27228
rect 8200 27172 8204 27228
rect 8140 27168 8204 27172
rect 14848 27228 14912 27232
rect 14848 27172 14852 27228
rect 14852 27172 14908 27228
rect 14908 27172 14912 27228
rect 14848 27168 14912 27172
rect 14928 27228 14992 27232
rect 14928 27172 14932 27228
rect 14932 27172 14988 27228
rect 14988 27172 14992 27228
rect 14928 27168 14992 27172
rect 15008 27228 15072 27232
rect 15008 27172 15012 27228
rect 15012 27172 15068 27228
rect 15068 27172 15072 27228
rect 15008 27168 15072 27172
rect 15088 27228 15152 27232
rect 15088 27172 15092 27228
rect 15092 27172 15148 27228
rect 15148 27172 15152 27228
rect 15088 27168 15152 27172
rect 21796 27228 21860 27232
rect 21796 27172 21800 27228
rect 21800 27172 21856 27228
rect 21856 27172 21860 27228
rect 21796 27168 21860 27172
rect 21876 27228 21940 27232
rect 21876 27172 21880 27228
rect 21880 27172 21936 27228
rect 21936 27172 21940 27228
rect 21876 27168 21940 27172
rect 21956 27228 22020 27232
rect 21956 27172 21960 27228
rect 21960 27172 22016 27228
rect 22016 27172 22020 27228
rect 21956 27168 22020 27172
rect 22036 27228 22100 27232
rect 22036 27172 22040 27228
rect 22040 27172 22096 27228
rect 22096 27172 22100 27228
rect 22036 27168 22100 27172
rect 4426 26684 4490 26688
rect 4426 26628 4430 26684
rect 4430 26628 4486 26684
rect 4486 26628 4490 26684
rect 4426 26624 4490 26628
rect 4506 26684 4570 26688
rect 4506 26628 4510 26684
rect 4510 26628 4566 26684
rect 4566 26628 4570 26684
rect 4506 26624 4570 26628
rect 4586 26684 4650 26688
rect 4586 26628 4590 26684
rect 4590 26628 4646 26684
rect 4646 26628 4650 26684
rect 4586 26624 4650 26628
rect 4666 26684 4730 26688
rect 4666 26628 4670 26684
rect 4670 26628 4726 26684
rect 4726 26628 4730 26684
rect 4666 26624 4730 26628
rect 11374 26684 11438 26688
rect 11374 26628 11378 26684
rect 11378 26628 11434 26684
rect 11434 26628 11438 26684
rect 11374 26624 11438 26628
rect 11454 26684 11518 26688
rect 11454 26628 11458 26684
rect 11458 26628 11514 26684
rect 11514 26628 11518 26684
rect 11454 26624 11518 26628
rect 11534 26684 11598 26688
rect 11534 26628 11538 26684
rect 11538 26628 11594 26684
rect 11594 26628 11598 26684
rect 11534 26624 11598 26628
rect 11614 26684 11678 26688
rect 11614 26628 11618 26684
rect 11618 26628 11674 26684
rect 11674 26628 11678 26684
rect 11614 26624 11678 26628
rect 18322 26684 18386 26688
rect 18322 26628 18326 26684
rect 18326 26628 18382 26684
rect 18382 26628 18386 26684
rect 18322 26624 18386 26628
rect 18402 26684 18466 26688
rect 18402 26628 18406 26684
rect 18406 26628 18462 26684
rect 18462 26628 18466 26684
rect 18402 26624 18466 26628
rect 18482 26684 18546 26688
rect 18482 26628 18486 26684
rect 18486 26628 18542 26684
rect 18542 26628 18546 26684
rect 18482 26624 18546 26628
rect 18562 26684 18626 26688
rect 18562 26628 18566 26684
rect 18566 26628 18622 26684
rect 18622 26628 18626 26684
rect 18562 26624 18626 26628
rect 25270 26684 25334 26688
rect 25270 26628 25274 26684
rect 25274 26628 25330 26684
rect 25330 26628 25334 26684
rect 25270 26624 25334 26628
rect 25350 26684 25414 26688
rect 25350 26628 25354 26684
rect 25354 26628 25410 26684
rect 25410 26628 25414 26684
rect 25350 26624 25414 26628
rect 25430 26684 25494 26688
rect 25430 26628 25434 26684
rect 25434 26628 25490 26684
rect 25490 26628 25494 26684
rect 25430 26624 25494 26628
rect 25510 26684 25574 26688
rect 25510 26628 25514 26684
rect 25514 26628 25570 26684
rect 25570 26628 25574 26684
rect 25510 26624 25574 26628
rect 7900 26140 7964 26144
rect 7900 26084 7904 26140
rect 7904 26084 7960 26140
rect 7960 26084 7964 26140
rect 7900 26080 7964 26084
rect 7980 26140 8044 26144
rect 7980 26084 7984 26140
rect 7984 26084 8040 26140
rect 8040 26084 8044 26140
rect 7980 26080 8044 26084
rect 8060 26140 8124 26144
rect 8060 26084 8064 26140
rect 8064 26084 8120 26140
rect 8120 26084 8124 26140
rect 8060 26080 8124 26084
rect 8140 26140 8204 26144
rect 8140 26084 8144 26140
rect 8144 26084 8200 26140
rect 8200 26084 8204 26140
rect 8140 26080 8204 26084
rect 14848 26140 14912 26144
rect 14848 26084 14852 26140
rect 14852 26084 14908 26140
rect 14908 26084 14912 26140
rect 14848 26080 14912 26084
rect 14928 26140 14992 26144
rect 14928 26084 14932 26140
rect 14932 26084 14988 26140
rect 14988 26084 14992 26140
rect 14928 26080 14992 26084
rect 15008 26140 15072 26144
rect 15008 26084 15012 26140
rect 15012 26084 15068 26140
rect 15068 26084 15072 26140
rect 15008 26080 15072 26084
rect 15088 26140 15152 26144
rect 15088 26084 15092 26140
rect 15092 26084 15148 26140
rect 15148 26084 15152 26140
rect 15088 26080 15152 26084
rect 21796 26140 21860 26144
rect 21796 26084 21800 26140
rect 21800 26084 21856 26140
rect 21856 26084 21860 26140
rect 21796 26080 21860 26084
rect 21876 26140 21940 26144
rect 21876 26084 21880 26140
rect 21880 26084 21936 26140
rect 21936 26084 21940 26140
rect 21876 26080 21940 26084
rect 21956 26140 22020 26144
rect 21956 26084 21960 26140
rect 21960 26084 22016 26140
rect 22016 26084 22020 26140
rect 21956 26080 22020 26084
rect 22036 26140 22100 26144
rect 22036 26084 22040 26140
rect 22040 26084 22096 26140
rect 22096 26084 22100 26140
rect 22036 26080 22100 26084
rect 4426 25596 4490 25600
rect 4426 25540 4430 25596
rect 4430 25540 4486 25596
rect 4486 25540 4490 25596
rect 4426 25536 4490 25540
rect 4506 25596 4570 25600
rect 4506 25540 4510 25596
rect 4510 25540 4566 25596
rect 4566 25540 4570 25596
rect 4506 25536 4570 25540
rect 4586 25596 4650 25600
rect 4586 25540 4590 25596
rect 4590 25540 4646 25596
rect 4646 25540 4650 25596
rect 4586 25536 4650 25540
rect 4666 25596 4730 25600
rect 4666 25540 4670 25596
rect 4670 25540 4726 25596
rect 4726 25540 4730 25596
rect 4666 25536 4730 25540
rect 11374 25596 11438 25600
rect 11374 25540 11378 25596
rect 11378 25540 11434 25596
rect 11434 25540 11438 25596
rect 11374 25536 11438 25540
rect 11454 25596 11518 25600
rect 11454 25540 11458 25596
rect 11458 25540 11514 25596
rect 11514 25540 11518 25596
rect 11454 25536 11518 25540
rect 11534 25596 11598 25600
rect 11534 25540 11538 25596
rect 11538 25540 11594 25596
rect 11594 25540 11598 25596
rect 11534 25536 11598 25540
rect 11614 25596 11678 25600
rect 11614 25540 11618 25596
rect 11618 25540 11674 25596
rect 11674 25540 11678 25596
rect 11614 25536 11678 25540
rect 18322 25596 18386 25600
rect 18322 25540 18326 25596
rect 18326 25540 18382 25596
rect 18382 25540 18386 25596
rect 18322 25536 18386 25540
rect 18402 25596 18466 25600
rect 18402 25540 18406 25596
rect 18406 25540 18462 25596
rect 18462 25540 18466 25596
rect 18402 25536 18466 25540
rect 18482 25596 18546 25600
rect 18482 25540 18486 25596
rect 18486 25540 18542 25596
rect 18542 25540 18546 25596
rect 18482 25536 18546 25540
rect 18562 25596 18626 25600
rect 18562 25540 18566 25596
rect 18566 25540 18622 25596
rect 18622 25540 18626 25596
rect 18562 25536 18626 25540
rect 25270 25596 25334 25600
rect 25270 25540 25274 25596
rect 25274 25540 25330 25596
rect 25330 25540 25334 25596
rect 25270 25536 25334 25540
rect 25350 25596 25414 25600
rect 25350 25540 25354 25596
rect 25354 25540 25410 25596
rect 25410 25540 25414 25596
rect 25350 25536 25414 25540
rect 25430 25596 25494 25600
rect 25430 25540 25434 25596
rect 25434 25540 25490 25596
rect 25490 25540 25494 25596
rect 25430 25536 25494 25540
rect 25510 25596 25574 25600
rect 25510 25540 25514 25596
rect 25514 25540 25570 25596
rect 25570 25540 25574 25596
rect 25510 25536 25574 25540
rect 7900 25052 7964 25056
rect 7900 24996 7904 25052
rect 7904 24996 7960 25052
rect 7960 24996 7964 25052
rect 7900 24992 7964 24996
rect 7980 25052 8044 25056
rect 7980 24996 7984 25052
rect 7984 24996 8040 25052
rect 8040 24996 8044 25052
rect 7980 24992 8044 24996
rect 8060 25052 8124 25056
rect 8060 24996 8064 25052
rect 8064 24996 8120 25052
rect 8120 24996 8124 25052
rect 8060 24992 8124 24996
rect 8140 25052 8204 25056
rect 8140 24996 8144 25052
rect 8144 24996 8200 25052
rect 8200 24996 8204 25052
rect 8140 24992 8204 24996
rect 14848 25052 14912 25056
rect 14848 24996 14852 25052
rect 14852 24996 14908 25052
rect 14908 24996 14912 25052
rect 14848 24992 14912 24996
rect 14928 25052 14992 25056
rect 14928 24996 14932 25052
rect 14932 24996 14988 25052
rect 14988 24996 14992 25052
rect 14928 24992 14992 24996
rect 15008 25052 15072 25056
rect 15008 24996 15012 25052
rect 15012 24996 15068 25052
rect 15068 24996 15072 25052
rect 15008 24992 15072 24996
rect 15088 25052 15152 25056
rect 15088 24996 15092 25052
rect 15092 24996 15148 25052
rect 15148 24996 15152 25052
rect 15088 24992 15152 24996
rect 21796 25052 21860 25056
rect 21796 24996 21800 25052
rect 21800 24996 21856 25052
rect 21856 24996 21860 25052
rect 21796 24992 21860 24996
rect 21876 25052 21940 25056
rect 21876 24996 21880 25052
rect 21880 24996 21936 25052
rect 21936 24996 21940 25052
rect 21876 24992 21940 24996
rect 21956 25052 22020 25056
rect 21956 24996 21960 25052
rect 21960 24996 22016 25052
rect 22016 24996 22020 25052
rect 21956 24992 22020 24996
rect 22036 25052 22100 25056
rect 22036 24996 22040 25052
rect 22040 24996 22096 25052
rect 22096 24996 22100 25052
rect 22036 24992 22100 24996
rect 4426 24508 4490 24512
rect 4426 24452 4430 24508
rect 4430 24452 4486 24508
rect 4486 24452 4490 24508
rect 4426 24448 4490 24452
rect 4506 24508 4570 24512
rect 4506 24452 4510 24508
rect 4510 24452 4566 24508
rect 4566 24452 4570 24508
rect 4506 24448 4570 24452
rect 4586 24508 4650 24512
rect 4586 24452 4590 24508
rect 4590 24452 4646 24508
rect 4646 24452 4650 24508
rect 4586 24448 4650 24452
rect 4666 24508 4730 24512
rect 4666 24452 4670 24508
rect 4670 24452 4726 24508
rect 4726 24452 4730 24508
rect 4666 24448 4730 24452
rect 11374 24508 11438 24512
rect 11374 24452 11378 24508
rect 11378 24452 11434 24508
rect 11434 24452 11438 24508
rect 11374 24448 11438 24452
rect 11454 24508 11518 24512
rect 11454 24452 11458 24508
rect 11458 24452 11514 24508
rect 11514 24452 11518 24508
rect 11454 24448 11518 24452
rect 11534 24508 11598 24512
rect 11534 24452 11538 24508
rect 11538 24452 11594 24508
rect 11594 24452 11598 24508
rect 11534 24448 11598 24452
rect 11614 24508 11678 24512
rect 11614 24452 11618 24508
rect 11618 24452 11674 24508
rect 11674 24452 11678 24508
rect 11614 24448 11678 24452
rect 18322 24508 18386 24512
rect 18322 24452 18326 24508
rect 18326 24452 18382 24508
rect 18382 24452 18386 24508
rect 18322 24448 18386 24452
rect 18402 24508 18466 24512
rect 18402 24452 18406 24508
rect 18406 24452 18462 24508
rect 18462 24452 18466 24508
rect 18402 24448 18466 24452
rect 18482 24508 18546 24512
rect 18482 24452 18486 24508
rect 18486 24452 18542 24508
rect 18542 24452 18546 24508
rect 18482 24448 18546 24452
rect 18562 24508 18626 24512
rect 18562 24452 18566 24508
rect 18566 24452 18622 24508
rect 18622 24452 18626 24508
rect 18562 24448 18626 24452
rect 25270 24508 25334 24512
rect 25270 24452 25274 24508
rect 25274 24452 25330 24508
rect 25330 24452 25334 24508
rect 25270 24448 25334 24452
rect 25350 24508 25414 24512
rect 25350 24452 25354 24508
rect 25354 24452 25410 24508
rect 25410 24452 25414 24508
rect 25350 24448 25414 24452
rect 25430 24508 25494 24512
rect 25430 24452 25434 24508
rect 25434 24452 25490 24508
rect 25490 24452 25494 24508
rect 25430 24448 25494 24452
rect 25510 24508 25574 24512
rect 25510 24452 25514 24508
rect 25514 24452 25570 24508
rect 25570 24452 25574 24508
rect 25510 24448 25574 24452
rect 7900 23964 7964 23968
rect 7900 23908 7904 23964
rect 7904 23908 7960 23964
rect 7960 23908 7964 23964
rect 7900 23904 7964 23908
rect 7980 23964 8044 23968
rect 7980 23908 7984 23964
rect 7984 23908 8040 23964
rect 8040 23908 8044 23964
rect 7980 23904 8044 23908
rect 8060 23964 8124 23968
rect 8060 23908 8064 23964
rect 8064 23908 8120 23964
rect 8120 23908 8124 23964
rect 8060 23904 8124 23908
rect 8140 23964 8204 23968
rect 8140 23908 8144 23964
rect 8144 23908 8200 23964
rect 8200 23908 8204 23964
rect 8140 23904 8204 23908
rect 14848 23964 14912 23968
rect 14848 23908 14852 23964
rect 14852 23908 14908 23964
rect 14908 23908 14912 23964
rect 14848 23904 14912 23908
rect 14928 23964 14992 23968
rect 14928 23908 14932 23964
rect 14932 23908 14988 23964
rect 14988 23908 14992 23964
rect 14928 23904 14992 23908
rect 15008 23964 15072 23968
rect 15008 23908 15012 23964
rect 15012 23908 15068 23964
rect 15068 23908 15072 23964
rect 15008 23904 15072 23908
rect 15088 23964 15152 23968
rect 15088 23908 15092 23964
rect 15092 23908 15148 23964
rect 15148 23908 15152 23964
rect 15088 23904 15152 23908
rect 21796 23964 21860 23968
rect 21796 23908 21800 23964
rect 21800 23908 21856 23964
rect 21856 23908 21860 23964
rect 21796 23904 21860 23908
rect 21876 23964 21940 23968
rect 21876 23908 21880 23964
rect 21880 23908 21936 23964
rect 21936 23908 21940 23964
rect 21876 23904 21940 23908
rect 21956 23964 22020 23968
rect 21956 23908 21960 23964
rect 21960 23908 22016 23964
rect 22016 23908 22020 23964
rect 21956 23904 22020 23908
rect 22036 23964 22100 23968
rect 22036 23908 22040 23964
rect 22040 23908 22096 23964
rect 22096 23908 22100 23964
rect 22036 23904 22100 23908
rect 4426 23420 4490 23424
rect 4426 23364 4430 23420
rect 4430 23364 4486 23420
rect 4486 23364 4490 23420
rect 4426 23360 4490 23364
rect 4506 23420 4570 23424
rect 4506 23364 4510 23420
rect 4510 23364 4566 23420
rect 4566 23364 4570 23420
rect 4506 23360 4570 23364
rect 4586 23420 4650 23424
rect 4586 23364 4590 23420
rect 4590 23364 4646 23420
rect 4646 23364 4650 23420
rect 4586 23360 4650 23364
rect 4666 23420 4730 23424
rect 4666 23364 4670 23420
rect 4670 23364 4726 23420
rect 4726 23364 4730 23420
rect 4666 23360 4730 23364
rect 11374 23420 11438 23424
rect 11374 23364 11378 23420
rect 11378 23364 11434 23420
rect 11434 23364 11438 23420
rect 11374 23360 11438 23364
rect 11454 23420 11518 23424
rect 11454 23364 11458 23420
rect 11458 23364 11514 23420
rect 11514 23364 11518 23420
rect 11454 23360 11518 23364
rect 11534 23420 11598 23424
rect 11534 23364 11538 23420
rect 11538 23364 11594 23420
rect 11594 23364 11598 23420
rect 11534 23360 11598 23364
rect 11614 23420 11678 23424
rect 11614 23364 11618 23420
rect 11618 23364 11674 23420
rect 11674 23364 11678 23420
rect 11614 23360 11678 23364
rect 18322 23420 18386 23424
rect 18322 23364 18326 23420
rect 18326 23364 18382 23420
rect 18382 23364 18386 23420
rect 18322 23360 18386 23364
rect 18402 23420 18466 23424
rect 18402 23364 18406 23420
rect 18406 23364 18462 23420
rect 18462 23364 18466 23420
rect 18402 23360 18466 23364
rect 18482 23420 18546 23424
rect 18482 23364 18486 23420
rect 18486 23364 18542 23420
rect 18542 23364 18546 23420
rect 18482 23360 18546 23364
rect 18562 23420 18626 23424
rect 18562 23364 18566 23420
rect 18566 23364 18622 23420
rect 18622 23364 18626 23420
rect 18562 23360 18626 23364
rect 25270 23420 25334 23424
rect 25270 23364 25274 23420
rect 25274 23364 25330 23420
rect 25330 23364 25334 23420
rect 25270 23360 25334 23364
rect 25350 23420 25414 23424
rect 25350 23364 25354 23420
rect 25354 23364 25410 23420
rect 25410 23364 25414 23420
rect 25350 23360 25414 23364
rect 25430 23420 25494 23424
rect 25430 23364 25434 23420
rect 25434 23364 25490 23420
rect 25490 23364 25494 23420
rect 25430 23360 25494 23364
rect 25510 23420 25574 23424
rect 25510 23364 25514 23420
rect 25514 23364 25570 23420
rect 25570 23364 25574 23420
rect 25510 23360 25574 23364
rect 7900 22876 7964 22880
rect 7900 22820 7904 22876
rect 7904 22820 7960 22876
rect 7960 22820 7964 22876
rect 7900 22816 7964 22820
rect 7980 22876 8044 22880
rect 7980 22820 7984 22876
rect 7984 22820 8040 22876
rect 8040 22820 8044 22876
rect 7980 22816 8044 22820
rect 8060 22876 8124 22880
rect 8060 22820 8064 22876
rect 8064 22820 8120 22876
rect 8120 22820 8124 22876
rect 8060 22816 8124 22820
rect 8140 22876 8204 22880
rect 8140 22820 8144 22876
rect 8144 22820 8200 22876
rect 8200 22820 8204 22876
rect 8140 22816 8204 22820
rect 14848 22876 14912 22880
rect 14848 22820 14852 22876
rect 14852 22820 14908 22876
rect 14908 22820 14912 22876
rect 14848 22816 14912 22820
rect 14928 22876 14992 22880
rect 14928 22820 14932 22876
rect 14932 22820 14988 22876
rect 14988 22820 14992 22876
rect 14928 22816 14992 22820
rect 15008 22876 15072 22880
rect 15008 22820 15012 22876
rect 15012 22820 15068 22876
rect 15068 22820 15072 22876
rect 15008 22816 15072 22820
rect 15088 22876 15152 22880
rect 15088 22820 15092 22876
rect 15092 22820 15148 22876
rect 15148 22820 15152 22876
rect 15088 22816 15152 22820
rect 21796 22876 21860 22880
rect 21796 22820 21800 22876
rect 21800 22820 21856 22876
rect 21856 22820 21860 22876
rect 21796 22816 21860 22820
rect 21876 22876 21940 22880
rect 21876 22820 21880 22876
rect 21880 22820 21936 22876
rect 21936 22820 21940 22876
rect 21876 22816 21940 22820
rect 21956 22876 22020 22880
rect 21956 22820 21960 22876
rect 21960 22820 22016 22876
rect 22016 22820 22020 22876
rect 21956 22816 22020 22820
rect 22036 22876 22100 22880
rect 22036 22820 22040 22876
rect 22040 22820 22096 22876
rect 22096 22820 22100 22876
rect 22036 22816 22100 22820
rect 4426 22332 4490 22336
rect 4426 22276 4430 22332
rect 4430 22276 4486 22332
rect 4486 22276 4490 22332
rect 4426 22272 4490 22276
rect 4506 22332 4570 22336
rect 4506 22276 4510 22332
rect 4510 22276 4566 22332
rect 4566 22276 4570 22332
rect 4506 22272 4570 22276
rect 4586 22332 4650 22336
rect 4586 22276 4590 22332
rect 4590 22276 4646 22332
rect 4646 22276 4650 22332
rect 4586 22272 4650 22276
rect 4666 22332 4730 22336
rect 4666 22276 4670 22332
rect 4670 22276 4726 22332
rect 4726 22276 4730 22332
rect 4666 22272 4730 22276
rect 11374 22332 11438 22336
rect 11374 22276 11378 22332
rect 11378 22276 11434 22332
rect 11434 22276 11438 22332
rect 11374 22272 11438 22276
rect 11454 22332 11518 22336
rect 11454 22276 11458 22332
rect 11458 22276 11514 22332
rect 11514 22276 11518 22332
rect 11454 22272 11518 22276
rect 11534 22332 11598 22336
rect 11534 22276 11538 22332
rect 11538 22276 11594 22332
rect 11594 22276 11598 22332
rect 11534 22272 11598 22276
rect 11614 22332 11678 22336
rect 11614 22276 11618 22332
rect 11618 22276 11674 22332
rect 11674 22276 11678 22332
rect 11614 22272 11678 22276
rect 18322 22332 18386 22336
rect 18322 22276 18326 22332
rect 18326 22276 18382 22332
rect 18382 22276 18386 22332
rect 18322 22272 18386 22276
rect 18402 22332 18466 22336
rect 18402 22276 18406 22332
rect 18406 22276 18462 22332
rect 18462 22276 18466 22332
rect 18402 22272 18466 22276
rect 18482 22332 18546 22336
rect 18482 22276 18486 22332
rect 18486 22276 18542 22332
rect 18542 22276 18546 22332
rect 18482 22272 18546 22276
rect 18562 22332 18626 22336
rect 18562 22276 18566 22332
rect 18566 22276 18622 22332
rect 18622 22276 18626 22332
rect 18562 22272 18626 22276
rect 25270 22332 25334 22336
rect 25270 22276 25274 22332
rect 25274 22276 25330 22332
rect 25330 22276 25334 22332
rect 25270 22272 25334 22276
rect 25350 22332 25414 22336
rect 25350 22276 25354 22332
rect 25354 22276 25410 22332
rect 25410 22276 25414 22332
rect 25350 22272 25414 22276
rect 25430 22332 25494 22336
rect 25430 22276 25434 22332
rect 25434 22276 25490 22332
rect 25490 22276 25494 22332
rect 25430 22272 25494 22276
rect 25510 22332 25574 22336
rect 25510 22276 25514 22332
rect 25514 22276 25570 22332
rect 25570 22276 25574 22332
rect 25510 22272 25574 22276
rect 7900 21788 7964 21792
rect 7900 21732 7904 21788
rect 7904 21732 7960 21788
rect 7960 21732 7964 21788
rect 7900 21728 7964 21732
rect 7980 21788 8044 21792
rect 7980 21732 7984 21788
rect 7984 21732 8040 21788
rect 8040 21732 8044 21788
rect 7980 21728 8044 21732
rect 8060 21788 8124 21792
rect 8060 21732 8064 21788
rect 8064 21732 8120 21788
rect 8120 21732 8124 21788
rect 8060 21728 8124 21732
rect 8140 21788 8204 21792
rect 8140 21732 8144 21788
rect 8144 21732 8200 21788
rect 8200 21732 8204 21788
rect 8140 21728 8204 21732
rect 14848 21788 14912 21792
rect 14848 21732 14852 21788
rect 14852 21732 14908 21788
rect 14908 21732 14912 21788
rect 14848 21728 14912 21732
rect 14928 21788 14992 21792
rect 14928 21732 14932 21788
rect 14932 21732 14988 21788
rect 14988 21732 14992 21788
rect 14928 21728 14992 21732
rect 15008 21788 15072 21792
rect 15008 21732 15012 21788
rect 15012 21732 15068 21788
rect 15068 21732 15072 21788
rect 15008 21728 15072 21732
rect 15088 21788 15152 21792
rect 15088 21732 15092 21788
rect 15092 21732 15148 21788
rect 15148 21732 15152 21788
rect 15088 21728 15152 21732
rect 21796 21788 21860 21792
rect 21796 21732 21800 21788
rect 21800 21732 21856 21788
rect 21856 21732 21860 21788
rect 21796 21728 21860 21732
rect 21876 21788 21940 21792
rect 21876 21732 21880 21788
rect 21880 21732 21936 21788
rect 21936 21732 21940 21788
rect 21876 21728 21940 21732
rect 21956 21788 22020 21792
rect 21956 21732 21960 21788
rect 21960 21732 22016 21788
rect 22016 21732 22020 21788
rect 21956 21728 22020 21732
rect 22036 21788 22100 21792
rect 22036 21732 22040 21788
rect 22040 21732 22096 21788
rect 22096 21732 22100 21788
rect 22036 21728 22100 21732
rect 4426 21244 4490 21248
rect 4426 21188 4430 21244
rect 4430 21188 4486 21244
rect 4486 21188 4490 21244
rect 4426 21184 4490 21188
rect 4506 21244 4570 21248
rect 4506 21188 4510 21244
rect 4510 21188 4566 21244
rect 4566 21188 4570 21244
rect 4506 21184 4570 21188
rect 4586 21244 4650 21248
rect 4586 21188 4590 21244
rect 4590 21188 4646 21244
rect 4646 21188 4650 21244
rect 4586 21184 4650 21188
rect 4666 21244 4730 21248
rect 4666 21188 4670 21244
rect 4670 21188 4726 21244
rect 4726 21188 4730 21244
rect 4666 21184 4730 21188
rect 11374 21244 11438 21248
rect 11374 21188 11378 21244
rect 11378 21188 11434 21244
rect 11434 21188 11438 21244
rect 11374 21184 11438 21188
rect 11454 21244 11518 21248
rect 11454 21188 11458 21244
rect 11458 21188 11514 21244
rect 11514 21188 11518 21244
rect 11454 21184 11518 21188
rect 11534 21244 11598 21248
rect 11534 21188 11538 21244
rect 11538 21188 11594 21244
rect 11594 21188 11598 21244
rect 11534 21184 11598 21188
rect 11614 21244 11678 21248
rect 11614 21188 11618 21244
rect 11618 21188 11674 21244
rect 11674 21188 11678 21244
rect 11614 21184 11678 21188
rect 18322 21244 18386 21248
rect 18322 21188 18326 21244
rect 18326 21188 18382 21244
rect 18382 21188 18386 21244
rect 18322 21184 18386 21188
rect 18402 21244 18466 21248
rect 18402 21188 18406 21244
rect 18406 21188 18462 21244
rect 18462 21188 18466 21244
rect 18402 21184 18466 21188
rect 18482 21244 18546 21248
rect 18482 21188 18486 21244
rect 18486 21188 18542 21244
rect 18542 21188 18546 21244
rect 18482 21184 18546 21188
rect 18562 21244 18626 21248
rect 18562 21188 18566 21244
rect 18566 21188 18622 21244
rect 18622 21188 18626 21244
rect 18562 21184 18626 21188
rect 25270 21244 25334 21248
rect 25270 21188 25274 21244
rect 25274 21188 25330 21244
rect 25330 21188 25334 21244
rect 25270 21184 25334 21188
rect 25350 21244 25414 21248
rect 25350 21188 25354 21244
rect 25354 21188 25410 21244
rect 25410 21188 25414 21244
rect 25350 21184 25414 21188
rect 25430 21244 25494 21248
rect 25430 21188 25434 21244
rect 25434 21188 25490 21244
rect 25490 21188 25494 21244
rect 25430 21184 25494 21188
rect 25510 21244 25574 21248
rect 25510 21188 25514 21244
rect 25514 21188 25570 21244
rect 25570 21188 25574 21244
rect 25510 21184 25574 21188
rect 7900 20700 7964 20704
rect 7900 20644 7904 20700
rect 7904 20644 7960 20700
rect 7960 20644 7964 20700
rect 7900 20640 7964 20644
rect 7980 20700 8044 20704
rect 7980 20644 7984 20700
rect 7984 20644 8040 20700
rect 8040 20644 8044 20700
rect 7980 20640 8044 20644
rect 8060 20700 8124 20704
rect 8060 20644 8064 20700
rect 8064 20644 8120 20700
rect 8120 20644 8124 20700
rect 8060 20640 8124 20644
rect 8140 20700 8204 20704
rect 8140 20644 8144 20700
rect 8144 20644 8200 20700
rect 8200 20644 8204 20700
rect 8140 20640 8204 20644
rect 14848 20700 14912 20704
rect 14848 20644 14852 20700
rect 14852 20644 14908 20700
rect 14908 20644 14912 20700
rect 14848 20640 14912 20644
rect 14928 20700 14992 20704
rect 14928 20644 14932 20700
rect 14932 20644 14988 20700
rect 14988 20644 14992 20700
rect 14928 20640 14992 20644
rect 15008 20700 15072 20704
rect 15008 20644 15012 20700
rect 15012 20644 15068 20700
rect 15068 20644 15072 20700
rect 15008 20640 15072 20644
rect 15088 20700 15152 20704
rect 15088 20644 15092 20700
rect 15092 20644 15148 20700
rect 15148 20644 15152 20700
rect 15088 20640 15152 20644
rect 21796 20700 21860 20704
rect 21796 20644 21800 20700
rect 21800 20644 21856 20700
rect 21856 20644 21860 20700
rect 21796 20640 21860 20644
rect 21876 20700 21940 20704
rect 21876 20644 21880 20700
rect 21880 20644 21936 20700
rect 21936 20644 21940 20700
rect 21876 20640 21940 20644
rect 21956 20700 22020 20704
rect 21956 20644 21960 20700
rect 21960 20644 22016 20700
rect 22016 20644 22020 20700
rect 21956 20640 22020 20644
rect 22036 20700 22100 20704
rect 22036 20644 22040 20700
rect 22040 20644 22096 20700
rect 22096 20644 22100 20700
rect 22036 20640 22100 20644
rect 4426 20156 4490 20160
rect 4426 20100 4430 20156
rect 4430 20100 4486 20156
rect 4486 20100 4490 20156
rect 4426 20096 4490 20100
rect 4506 20156 4570 20160
rect 4506 20100 4510 20156
rect 4510 20100 4566 20156
rect 4566 20100 4570 20156
rect 4506 20096 4570 20100
rect 4586 20156 4650 20160
rect 4586 20100 4590 20156
rect 4590 20100 4646 20156
rect 4646 20100 4650 20156
rect 4586 20096 4650 20100
rect 4666 20156 4730 20160
rect 4666 20100 4670 20156
rect 4670 20100 4726 20156
rect 4726 20100 4730 20156
rect 4666 20096 4730 20100
rect 11374 20156 11438 20160
rect 11374 20100 11378 20156
rect 11378 20100 11434 20156
rect 11434 20100 11438 20156
rect 11374 20096 11438 20100
rect 11454 20156 11518 20160
rect 11454 20100 11458 20156
rect 11458 20100 11514 20156
rect 11514 20100 11518 20156
rect 11454 20096 11518 20100
rect 11534 20156 11598 20160
rect 11534 20100 11538 20156
rect 11538 20100 11594 20156
rect 11594 20100 11598 20156
rect 11534 20096 11598 20100
rect 11614 20156 11678 20160
rect 11614 20100 11618 20156
rect 11618 20100 11674 20156
rect 11674 20100 11678 20156
rect 11614 20096 11678 20100
rect 18322 20156 18386 20160
rect 18322 20100 18326 20156
rect 18326 20100 18382 20156
rect 18382 20100 18386 20156
rect 18322 20096 18386 20100
rect 18402 20156 18466 20160
rect 18402 20100 18406 20156
rect 18406 20100 18462 20156
rect 18462 20100 18466 20156
rect 18402 20096 18466 20100
rect 18482 20156 18546 20160
rect 18482 20100 18486 20156
rect 18486 20100 18542 20156
rect 18542 20100 18546 20156
rect 18482 20096 18546 20100
rect 18562 20156 18626 20160
rect 18562 20100 18566 20156
rect 18566 20100 18622 20156
rect 18622 20100 18626 20156
rect 18562 20096 18626 20100
rect 25270 20156 25334 20160
rect 25270 20100 25274 20156
rect 25274 20100 25330 20156
rect 25330 20100 25334 20156
rect 25270 20096 25334 20100
rect 25350 20156 25414 20160
rect 25350 20100 25354 20156
rect 25354 20100 25410 20156
rect 25410 20100 25414 20156
rect 25350 20096 25414 20100
rect 25430 20156 25494 20160
rect 25430 20100 25434 20156
rect 25434 20100 25490 20156
rect 25490 20100 25494 20156
rect 25430 20096 25494 20100
rect 25510 20156 25574 20160
rect 25510 20100 25514 20156
rect 25514 20100 25570 20156
rect 25570 20100 25574 20156
rect 25510 20096 25574 20100
rect 7900 19612 7964 19616
rect 7900 19556 7904 19612
rect 7904 19556 7960 19612
rect 7960 19556 7964 19612
rect 7900 19552 7964 19556
rect 7980 19612 8044 19616
rect 7980 19556 7984 19612
rect 7984 19556 8040 19612
rect 8040 19556 8044 19612
rect 7980 19552 8044 19556
rect 8060 19612 8124 19616
rect 8060 19556 8064 19612
rect 8064 19556 8120 19612
rect 8120 19556 8124 19612
rect 8060 19552 8124 19556
rect 8140 19612 8204 19616
rect 8140 19556 8144 19612
rect 8144 19556 8200 19612
rect 8200 19556 8204 19612
rect 8140 19552 8204 19556
rect 14848 19612 14912 19616
rect 14848 19556 14852 19612
rect 14852 19556 14908 19612
rect 14908 19556 14912 19612
rect 14848 19552 14912 19556
rect 14928 19612 14992 19616
rect 14928 19556 14932 19612
rect 14932 19556 14988 19612
rect 14988 19556 14992 19612
rect 14928 19552 14992 19556
rect 15008 19612 15072 19616
rect 15008 19556 15012 19612
rect 15012 19556 15068 19612
rect 15068 19556 15072 19612
rect 15008 19552 15072 19556
rect 15088 19612 15152 19616
rect 15088 19556 15092 19612
rect 15092 19556 15148 19612
rect 15148 19556 15152 19612
rect 15088 19552 15152 19556
rect 21796 19612 21860 19616
rect 21796 19556 21800 19612
rect 21800 19556 21856 19612
rect 21856 19556 21860 19612
rect 21796 19552 21860 19556
rect 21876 19612 21940 19616
rect 21876 19556 21880 19612
rect 21880 19556 21936 19612
rect 21936 19556 21940 19612
rect 21876 19552 21940 19556
rect 21956 19612 22020 19616
rect 21956 19556 21960 19612
rect 21960 19556 22016 19612
rect 22016 19556 22020 19612
rect 21956 19552 22020 19556
rect 22036 19612 22100 19616
rect 22036 19556 22040 19612
rect 22040 19556 22096 19612
rect 22096 19556 22100 19612
rect 22036 19552 22100 19556
rect 4426 19068 4490 19072
rect 4426 19012 4430 19068
rect 4430 19012 4486 19068
rect 4486 19012 4490 19068
rect 4426 19008 4490 19012
rect 4506 19068 4570 19072
rect 4506 19012 4510 19068
rect 4510 19012 4566 19068
rect 4566 19012 4570 19068
rect 4506 19008 4570 19012
rect 4586 19068 4650 19072
rect 4586 19012 4590 19068
rect 4590 19012 4646 19068
rect 4646 19012 4650 19068
rect 4586 19008 4650 19012
rect 4666 19068 4730 19072
rect 4666 19012 4670 19068
rect 4670 19012 4726 19068
rect 4726 19012 4730 19068
rect 4666 19008 4730 19012
rect 11374 19068 11438 19072
rect 11374 19012 11378 19068
rect 11378 19012 11434 19068
rect 11434 19012 11438 19068
rect 11374 19008 11438 19012
rect 11454 19068 11518 19072
rect 11454 19012 11458 19068
rect 11458 19012 11514 19068
rect 11514 19012 11518 19068
rect 11454 19008 11518 19012
rect 11534 19068 11598 19072
rect 11534 19012 11538 19068
rect 11538 19012 11594 19068
rect 11594 19012 11598 19068
rect 11534 19008 11598 19012
rect 11614 19068 11678 19072
rect 11614 19012 11618 19068
rect 11618 19012 11674 19068
rect 11674 19012 11678 19068
rect 11614 19008 11678 19012
rect 18322 19068 18386 19072
rect 18322 19012 18326 19068
rect 18326 19012 18382 19068
rect 18382 19012 18386 19068
rect 18322 19008 18386 19012
rect 18402 19068 18466 19072
rect 18402 19012 18406 19068
rect 18406 19012 18462 19068
rect 18462 19012 18466 19068
rect 18402 19008 18466 19012
rect 18482 19068 18546 19072
rect 18482 19012 18486 19068
rect 18486 19012 18542 19068
rect 18542 19012 18546 19068
rect 18482 19008 18546 19012
rect 18562 19068 18626 19072
rect 18562 19012 18566 19068
rect 18566 19012 18622 19068
rect 18622 19012 18626 19068
rect 18562 19008 18626 19012
rect 25270 19068 25334 19072
rect 25270 19012 25274 19068
rect 25274 19012 25330 19068
rect 25330 19012 25334 19068
rect 25270 19008 25334 19012
rect 25350 19068 25414 19072
rect 25350 19012 25354 19068
rect 25354 19012 25410 19068
rect 25410 19012 25414 19068
rect 25350 19008 25414 19012
rect 25430 19068 25494 19072
rect 25430 19012 25434 19068
rect 25434 19012 25490 19068
rect 25490 19012 25494 19068
rect 25430 19008 25494 19012
rect 25510 19068 25574 19072
rect 25510 19012 25514 19068
rect 25514 19012 25570 19068
rect 25570 19012 25574 19068
rect 25510 19008 25574 19012
rect 7900 18524 7964 18528
rect 7900 18468 7904 18524
rect 7904 18468 7960 18524
rect 7960 18468 7964 18524
rect 7900 18464 7964 18468
rect 7980 18524 8044 18528
rect 7980 18468 7984 18524
rect 7984 18468 8040 18524
rect 8040 18468 8044 18524
rect 7980 18464 8044 18468
rect 8060 18524 8124 18528
rect 8060 18468 8064 18524
rect 8064 18468 8120 18524
rect 8120 18468 8124 18524
rect 8060 18464 8124 18468
rect 8140 18524 8204 18528
rect 8140 18468 8144 18524
rect 8144 18468 8200 18524
rect 8200 18468 8204 18524
rect 8140 18464 8204 18468
rect 14848 18524 14912 18528
rect 14848 18468 14852 18524
rect 14852 18468 14908 18524
rect 14908 18468 14912 18524
rect 14848 18464 14912 18468
rect 14928 18524 14992 18528
rect 14928 18468 14932 18524
rect 14932 18468 14988 18524
rect 14988 18468 14992 18524
rect 14928 18464 14992 18468
rect 15008 18524 15072 18528
rect 15008 18468 15012 18524
rect 15012 18468 15068 18524
rect 15068 18468 15072 18524
rect 15008 18464 15072 18468
rect 15088 18524 15152 18528
rect 15088 18468 15092 18524
rect 15092 18468 15148 18524
rect 15148 18468 15152 18524
rect 15088 18464 15152 18468
rect 21796 18524 21860 18528
rect 21796 18468 21800 18524
rect 21800 18468 21856 18524
rect 21856 18468 21860 18524
rect 21796 18464 21860 18468
rect 21876 18524 21940 18528
rect 21876 18468 21880 18524
rect 21880 18468 21936 18524
rect 21936 18468 21940 18524
rect 21876 18464 21940 18468
rect 21956 18524 22020 18528
rect 21956 18468 21960 18524
rect 21960 18468 22016 18524
rect 22016 18468 22020 18524
rect 21956 18464 22020 18468
rect 22036 18524 22100 18528
rect 22036 18468 22040 18524
rect 22040 18468 22096 18524
rect 22096 18468 22100 18524
rect 22036 18464 22100 18468
rect 4426 17980 4490 17984
rect 4426 17924 4430 17980
rect 4430 17924 4486 17980
rect 4486 17924 4490 17980
rect 4426 17920 4490 17924
rect 4506 17980 4570 17984
rect 4506 17924 4510 17980
rect 4510 17924 4566 17980
rect 4566 17924 4570 17980
rect 4506 17920 4570 17924
rect 4586 17980 4650 17984
rect 4586 17924 4590 17980
rect 4590 17924 4646 17980
rect 4646 17924 4650 17980
rect 4586 17920 4650 17924
rect 4666 17980 4730 17984
rect 4666 17924 4670 17980
rect 4670 17924 4726 17980
rect 4726 17924 4730 17980
rect 4666 17920 4730 17924
rect 11374 17980 11438 17984
rect 11374 17924 11378 17980
rect 11378 17924 11434 17980
rect 11434 17924 11438 17980
rect 11374 17920 11438 17924
rect 11454 17980 11518 17984
rect 11454 17924 11458 17980
rect 11458 17924 11514 17980
rect 11514 17924 11518 17980
rect 11454 17920 11518 17924
rect 11534 17980 11598 17984
rect 11534 17924 11538 17980
rect 11538 17924 11594 17980
rect 11594 17924 11598 17980
rect 11534 17920 11598 17924
rect 11614 17980 11678 17984
rect 11614 17924 11618 17980
rect 11618 17924 11674 17980
rect 11674 17924 11678 17980
rect 11614 17920 11678 17924
rect 18322 17980 18386 17984
rect 18322 17924 18326 17980
rect 18326 17924 18382 17980
rect 18382 17924 18386 17980
rect 18322 17920 18386 17924
rect 18402 17980 18466 17984
rect 18402 17924 18406 17980
rect 18406 17924 18462 17980
rect 18462 17924 18466 17980
rect 18402 17920 18466 17924
rect 18482 17980 18546 17984
rect 18482 17924 18486 17980
rect 18486 17924 18542 17980
rect 18542 17924 18546 17980
rect 18482 17920 18546 17924
rect 18562 17980 18626 17984
rect 18562 17924 18566 17980
rect 18566 17924 18622 17980
rect 18622 17924 18626 17980
rect 18562 17920 18626 17924
rect 25270 17980 25334 17984
rect 25270 17924 25274 17980
rect 25274 17924 25330 17980
rect 25330 17924 25334 17980
rect 25270 17920 25334 17924
rect 25350 17980 25414 17984
rect 25350 17924 25354 17980
rect 25354 17924 25410 17980
rect 25410 17924 25414 17980
rect 25350 17920 25414 17924
rect 25430 17980 25494 17984
rect 25430 17924 25434 17980
rect 25434 17924 25490 17980
rect 25490 17924 25494 17980
rect 25430 17920 25494 17924
rect 25510 17980 25574 17984
rect 25510 17924 25514 17980
rect 25514 17924 25570 17980
rect 25570 17924 25574 17980
rect 25510 17920 25574 17924
rect 7900 17436 7964 17440
rect 7900 17380 7904 17436
rect 7904 17380 7960 17436
rect 7960 17380 7964 17436
rect 7900 17376 7964 17380
rect 7980 17436 8044 17440
rect 7980 17380 7984 17436
rect 7984 17380 8040 17436
rect 8040 17380 8044 17436
rect 7980 17376 8044 17380
rect 8060 17436 8124 17440
rect 8060 17380 8064 17436
rect 8064 17380 8120 17436
rect 8120 17380 8124 17436
rect 8060 17376 8124 17380
rect 8140 17436 8204 17440
rect 8140 17380 8144 17436
rect 8144 17380 8200 17436
rect 8200 17380 8204 17436
rect 8140 17376 8204 17380
rect 14848 17436 14912 17440
rect 14848 17380 14852 17436
rect 14852 17380 14908 17436
rect 14908 17380 14912 17436
rect 14848 17376 14912 17380
rect 14928 17436 14992 17440
rect 14928 17380 14932 17436
rect 14932 17380 14988 17436
rect 14988 17380 14992 17436
rect 14928 17376 14992 17380
rect 15008 17436 15072 17440
rect 15008 17380 15012 17436
rect 15012 17380 15068 17436
rect 15068 17380 15072 17436
rect 15008 17376 15072 17380
rect 15088 17436 15152 17440
rect 15088 17380 15092 17436
rect 15092 17380 15148 17436
rect 15148 17380 15152 17436
rect 15088 17376 15152 17380
rect 21796 17436 21860 17440
rect 21796 17380 21800 17436
rect 21800 17380 21856 17436
rect 21856 17380 21860 17436
rect 21796 17376 21860 17380
rect 21876 17436 21940 17440
rect 21876 17380 21880 17436
rect 21880 17380 21936 17436
rect 21936 17380 21940 17436
rect 21876 17376 21940 17380
rect 21956 17436 22020 17440
rect 21956 17380 21960 17436
rect 21960 17380 22016 17436
rect 22016 17380 22020 17436
rect 21956 17376 22020 17380
rect 22036 17436 22100 17440
rect 22036 17380 22040 17436
rect 22040 17380 22096 17436
rect 22096 17380 22100 17436
rect 22036 17376 22100 17380
rect 4426 16892 4490 16896
rect 4426 16836 4430 16892
rect 4430 16836 4486 16892
rect 4486 16836 4490 16892
rect 4426 16832 4490 16836
rect 4506 16892 4570 16896
rect 4506 16836 4510 16892
rect 4510 16836 4566 16892
rect 4566 16836 4570 16892
rect 4506 16832 4570 16836
rect 4586 16892 4650 16896
rect 4586 16836 4590 16892
rect 4590 16836 4646 16892
rect 4646 16836 4650 16892
rect 4586 16832 4650 16836
rect 4666 16892 4730 16896
rect 4666 16836 4670 16892
rect 4670 16836 4726 16892
rect 4726 16836 4730 16892
rect 4666 16832 4730 16836
rect 11374 16892 11438 16896
rect 11374 16836 11378 16892
rect 11378 16836 11434 16892
rect 11434 16836 11438 16892
rect 11374 16832 11438 16836
rect 11454 16892 11518 16896
rect 11454 16836 11458 16892
rect 11458 16836 11514 16892
rect 11514 16836 11518 16892
rect 11454 16832 11518 16836
rect 11534 16892 11598 16896
rect 11534 16836 11538 16892
rect 11538 16836 11594 16892
rect 11594 16836 11598 16892
rect 11534 16832 11598 16836
rect 11614 16892 11678 16896
rect 11614 16836 11618 16892
rect 11618 16836 11674 16892
rect 11674 16836 11678 16892
rect 11614 16832 11678 16836
rect 18322 16892 18386 16896
rect 18322 16836 18326 16892
rect 18326 16836 18382 16892
rect 18382 16836 18386 16892
rect 18322 16832 18386 16836
rect 18402 16892 18466 16896
rect 18402 16836 18406 16892
rect 18406 16836 18462 16892
rect 18462 16836 18466 16892
rect 18402 16832 18466 16836
rect 18482 16892 18546 16896
rect 18482 16836 18486 16892
rect 18486 16836 18542 16892
rect 18542 16836 18546 16892
rect 18482 16832 18546 16836
rect 18562 16892 18626 16896
rect 18562 16836 18566 16892
rect 18566 16836 18622 16892
rect 18622 16836 18626 16892
rect 18562 16832 18626 16836
rect 25270 16892 25334 16896
rect 25270 16836 25274 16892
rect 25274 16836 25330 16892
rect 25330 16836 25334 16892
rect 25270 16832 25334 16836
rect 25350 16892 25414 16896
rect 25350 16836 25354 16892
rect 25354 16836 25410 16892
rect 25410 16836 25414 16892
rect 25350 16832 25414 16836
rect 25430 16892 25494 16896
rect 25430 16836 25434 16892
rect 25434 16836 25490 16892
rect 25490 16836 25494 16892
rect 25430 16832 25494 16836
rect 25510 16892 25574 16896
rect 25510 16836 25514 16892
rect 25514 16836 25570 16892
rect 25570 16836 25574 16892
rect 25510 16832 25574 16836
rect 7900 16348 7964 16352
rect 7900 16292 7904 16348
rect 7904 16292 7960 16348
rect 7960 16292 7964 16348
rect 7900 16288 7964 16292
rect 7980 16348 8044 16352
rect 7980 16292 7984 16348
rect 7984 16292 8040 16348
rect 8040 16292 8044 16348
rect 7980 16288 8044 16292
rect 8060 16348 8124 16352
rect 8060 16292 8064 16348
rect 8064 16292 8120 16348
rect 8120 16292 8124 16348
rect 8060 16288 8124 16292
rect 8140 16348 8204 16352
rect 8140 16292 8144 16348
rect 8144 16292 8200 16348
rect 8200 16292 8204 16348
rect 8140 16288 8204 16292
rect 14848 16348 14912 16352
rect 14848 16292 14852 16348
rect 14852 16292 14908 16348
rect 14908 16292 14912 16348
rect 14848 16288 14912 16292
rect 14928 16348 14992 16352
rect 14928 16292 14932 16348
rect 14932 16292 14988 16348
rect 14988 16292 14992 16348
rect 14928 16288 14992 16292
rect 15008 16348 15072 16352
rect 15008 16292 15012 16348
rect 15012 16292 15068 16348
rect 15068 16292 15072 16348
rect 15008 16288 15072 16292
rect 15088 16348 15152 16352
rect 15088 16292 15092 16348
rect 15092 16292 15148 16348
rect 15148 16292 15152 16348
rect 15088 16288 15152 16292
rect 21796 16348 21860 16352
rect 21796 16292 21800 16348
rect 21800 16292 21856 16348
rect 21856 16292 21860 16348
rect 21796 16288 21860 16292
rect 21876 16348 21940 16352
rect 21876 16292 21880 16348
rect 21880 16292 21936 16348
rect 21936 16292 21940 16348
rect 21876 16288 21940 16292
rect 21956 16348 22020 16352
rect 21956 16292 21960 16348
rect 21960 16292 22016 16348
rect 22016 16292 22020 16348
rect 21956 16288 22020 16292
rect 22036 16348 22100 16352
rect 22036 16292 22040 16348
rect 22040 16292 22096 16348
rect 22096 16292 22100 16348
rect 22036 16288 22100 16292
rect 4426 15804 4490 15808
rect 4426 15748 4430 15804
rect 4430 15748 4486 15804
rect 4486 15748 4490 15804
rect 4426 15744 4490 15748
rect 4506 15804 4570 15808
rect 4506 15748 4510 15804
rect 4510 15748 4566 15804
rect 4566 15748 4570 15804
rect 4506 15744 4570 15748
rect 4586 15804 4650 15808
rect 4586 15748 4590 15804
rect 4590 15748 4646 15804
rect 4646 15748 4650 15804
rect 4586 15744 4650 15748
rect 4666 15804 4730 15808
rect 4666 15748 4670 15804
rect 4670 15748 4726 15804
rect 4726 15748 4730 15804
rect 4666 15744 4730 15748
rect 11374 15804 11438 15808
rect 11374 15748 11378 15804
rect 11378 15748 11434 15804
rect 11434 15748 11438 15804
rect 11374 15744 11438 15748
rect 11454 15804 11518 15808
rect 11454 15748 11458 15804
rect 11458 15748 11514 15804
rect 11514 15748 11518 15804
rect 11454 15744 11518 15748
rect 11534 15804 11598 15808
rect 11534 15748 11538 15804
rect 11538 15748 11594 15804
rect 11594 15748 11598 15804
rect 11534 15744 11598 15748
rect 11614 15804 11678 15808
rect 11614 15748 11618 15804
rect 11618 15748 11674 15804
rect 11674 15748 11678 15804
rect 11614 15744 11678 15748
rect 18322 15804 18386 15808
rect 18322 15748 18326 15804
rect 18326 15748 18382 15804
rect 18382 15748 18386 15804
rect 18322 15744 18386 15748
rect 18402 15804 18466 15808
rect 18402 15748 18406 15804
rect 18406 15748 18462 15804
rect 18462 15748 18466 15804
rect 18402 15744 18466 15748
rect 18482 15804 18546 15808
rect 18482 15748 18486 15804
rect 18486 15748 18542 15804
rect 18542 15748 18546 15804
rect 18482 15744 18546 15748
rect 18562 15804 18626 15808
rect 18562 15748 18566 15804
rect 18566 15748 18622 15804
rect 18622 15748 18626 15804
rect 18562 15744 18626 15748
rect 25270 15804 25334 15808
rect 25270 15748 25274 15804
rect 25274 15748 25330 15804
rect 25330 15748 25334 15804
rect 25270 15744 25334 15748
rect 25350 15804 25414 15808
rect 25350 15748 25354 15804
rect 25354 15748 25410 15804
rect 25410 15748 25414 15804
rect 25350 15744 25414 15748
rect 25430 15804 25494 15808
rect 25430 15748 25434 15804
rect 25434 15748 25490 15804
rect 25490 15748 25494 15804
rect 25430 15744 25494 15748
rect 25510 15804 25574 15808
rect 25510 15748 25514 15804
rect 25514 15748 25570 15804
rect 25570 15748 25574 15804
rect 25510 15744 25574 15748
rect 7900 15260 7964 15264
rect 7900 15204 7904 15260
rect 7904 15204 7960 15260
rect 7960 15204 7964 15260
rect 7900 15200 7964 15204
rect 7980 15260 8044 15264
rect 7980 15204 7984 15260
rect 7984 15204 8040 15260
rect 8040 15204 8044 15260
rect 7980 15200 8044 15204
rect 8060 15260 8124 15264
rect 8060 15204 8064 15260
rect 8064 15204 8120 15260
rect 8120 15204 8124 15260
rect 8060 15200 8124 15204
rect 8140 15260 8204 15264
rect 8140 15204 8144 15260
rect 8144 15204 8200 15260
rect 8200 15204 8204 15260
rect 8140 15200 8204 15204
rect 14848 15260 14912 15264
rect 14848 15204 14852 15260
rect 14852 15204 14908 15260
rect 14908 15204 14912 15260
rect 14848 15200 14912 15204
rect 14928 15260 14992 15264
rect 14928 15204 14932 15260
rect 14932 15204 14988 15260
rect 14988 15204 14992 15260
rect 14928 15200 14992 15204
rect 15008 15260 15072 15264
rect 15008 15204 15012 15260
rect 15012 15204 15068 15260
rect 15068 15204 15072 15260
rect 15008 15200 15072 15204
rect 15088 15260 15152 15264
rect 15088 15204 15092 15260
rect 15092 15204 15148 15260
rect 15148 15204 15152 15260
rect 15088 15200 15152 15204
rect 21796 15260 21860 15264
rect 21796 15204 21800 15260
rect 21800 15204 21856 15260
rect 21856 15204 21860 15260
rect 21796 15200 21860 15204
rect 21876 15260 21940 15264
rect 21876 15204 21880 15260
rect 21880 15204 21936 15260
rect 21936 15204 21940 15260
rect 21876 15200 21940 15204
rect 21956 15260 22020 15264
rect 21956 15204 21960 15260
rect 21960 15204 22016 15260
rect 22016 15204 22020 15260
rect 21956 15200 22020 15204
rect 22036 15260 22100 15264
rect 22036 15204 22040 15260
rect 22040 15204 22096 15260
rect 22096 15204 22100 15260
rect 22036 15200 22100 15204
rect 4426 14716 4490 14720
rect 4426 14660 4430 14716
rect 4430 14660 4486 14716
rect 4486 14660 4490 14716
rect 4426 14656 4490 14660
rect 4506 14716 4570 14720
rect 4506 14660 4510 14716
rect 4510 14660 4566 14716
rect 4566 14660 4570 14716
rect 4506 14656 4570 14660
rect 4586 14716 4650 14720
rect 4586 14660 4590 14716
rect 4590 14660 4646 14716
rect 4646 14660 4650 14716
rect 4586 14656 4650 14660
rect 4666 14716 4730 14720
rect 4666 14660 4670 14716
rect 4670 14660 4726 14716
rect 4726 14660 4730 14716
rect 4666 14656 4730 14660
rect 11374 14716 11438 14720
rect 11374 14660 11378 14716
rect 11378 14660 11434 14716
rect 11434 14660 11438 14716
rect 11374 14656 11438 14660
rect 11454 14716 11518 14720
rect 11454 14660 11458 14716
rect 11458 14660 11514 14716
rect 11514 14660 11518 14716
rect 11454 14656 11518 14660
rect 11534 14716 11598 14720
rect 11534 14660 11538 14716
rect 11538 14660 11594 14716
rect 11594 14660 11598 14716
rect 11534 14656 11598 14660
rect 11614 14716 11678 14720
rect 11614 14660 11618 14716
rect 11618 14660 11674 14716
rect 11674 14660 11678 14716
rect 11614 14656 11678 14660
rect 18322 14716 18386 14720
rect 18322 14660 18326 14716
rect 18326 14660 18382 14716
rect 18382 14660 18386 14716
rect 18322 14656 18386 14660
rect 18402 14716 18466 14720
rect 18402 14660 18406 14716
rect 18406 14660 18462 14716
rect 18462 14660 18466 14716
rect 18402 14656 18466 14660
rect 18482 14716 18546 14720
rect 18482 14660 18486 14716
rect 18486 14660 18542 14716
rect 18542 14660 18546 14716
rect 18482 14656 18546 14660
rect 18562 14716 18626 14720
rect 18562 14660 18566 14716
rect 18566 14660 18622 14716
rect 18622 14660 18626 14716
rect 18562 14656 18626 14660
rect 25270 14716 25334 14720
rect 25270 14660 25274 14716
rect 25274 14660 25330 14716
rect 25330 14660 25334 14716
rect 25270 14656 25334 14660
rect 25350 14716 25414 14720
rect 25350 14660 25354 14716
rect 25354 14660 25410 14716
rect 25410 14660 25414 14716
rect 25350 14656 25414 14660
rect 25430 14716 25494 14720
rect 25430 14660 25434 14716
rect 25434 14660 25490 14716
rect 25490 14660 25494 14716
rect 25430 14656 25494 14660
rect 25510 14716 25574 14720
rect 25510 14660 25514 14716
rect 25514 14660 25570 14716
rect 25570 14660 25574 14716
rect 25510 14656 25574 14660
rect 7900 14172 7964 14176
rect 7900 14116 7904 14172
rect 7904 14116 7960 14172
rect 7960 14116 7964 14172
rect 7900 14112 7964 14116
rect 7980 14172 8044 14176
rect 7980 14116 7984 14172
rect 7984 14116 8040 14172
rect 8040 14116 8044 14172
rect 7980 14112 8044 14116
rect 8060 14172 8124 14176
rect 8060 14116 8064 14172
rect 8064 14116 8120 14172
rect 8120 14116 8124 14172
rect 8060 14112 8124 14116
rect 8140 14172 8204 14176
rect 8140 14116 8144 14172
rect 8144 14116 8200 14172
rect 8200 14116 8204 14172
rect 8140 14112 8204 14116
rect 14848 14172 14912 14176
rect 14848 14116 14852 14172
rect 14852 14116 14908 14172
rect 14908 14116 14912 14172
rect 14848 14112 14912 14116
rect 14928 14172 14992 14176
rect 14928 14116 14932 14172
rect 14932 14116 14988 14172
rect 14988 14116 14992 14172
rect 14928 14112 14992 14116
rect 15008 14172 15072 14176
rect 15008 14116 15012 14172
rect 15012 14116 15068 14172
rect 15068 14116 15072 14172
rect 15008 14112 15072 14116
rect 15088 14172 15152 14176
rect 15088 14116 15092 14172
rect 15092 14116 15148 14172
rect 15148 14116 15152 14172
rect 15088 14112 15152 14116
rect 21796 14172 21860 14176
rect 21796 14116 21800 14172
rect 21800 14116 21856 14172
rect 21856 14116 21860 14172
rect 21796 14112 21860 14116
rect 21876 14172 21940 14176
rect 21876 14116 21880 14172
rect 21880 14116 21936 14172
rect 21936 14116 21940 14172
rect 21876 14112 21940 14116
rect 21956 14172 22020 14176
rect 21956 14116 21960 14172
rect 21960 14116 22016 14172
rect 22016 14116 22020 14172
rect 21956 14112 22020 14116
rect 22036 14172 22100 14176
rect 22036 14116 22040 14172
rect 22040 14116 22096 14172
rect 22096 14116 22100 14172
rect 22036 14112 22100 14116
rect 4426 13628 4490 13632
rect 4426 13572 4430 13628
rect 4430 13572 4486 13628
rect 4486 13572 4490 13628
rect 4426 13568 4490 13572
rect 4506 13628 4570 13632
rect 4506 13572 4510 13628
rect 4510 13572 4566 13628
rect 4566 13572 4570 13628
rect 4506 13568 4570 13572
rect 4586 13628 4650 13632
rect 4586 13572 4590 13628
rect 4590 13572 4646 13628
rect 4646 13572 4650 13628
rect 4586 13568 4650 13572
rect 4666 13628 4730 13632
rect 4666 13572 4670 13628
rect 4670 13572 4726 13628
rect 4726 13572 4730 13628
rect 4666 13568 4730 13572
rect 11374 13628 11438 13632
rect 11374 13572 11378 13628
rect 11378 13572 11434 13628
rect 11434 13572 11438 13628
rect 11374 13568 11438 13572
rect 11454 13628 11518 13632
rect 11454 13572 11458 13628
rect 11458 13572 11514 13628
rect 11514 13572 11518 13628
rect 11454 13568 11518 13572
rect 11534 13628 11598 13632
rect 11534 13572 11538 13628
rect 11538 13572 11594 13628
rect 11594 13572 11598 13628
rect 11534 13568 11598 13572
rect 11614 13628 11678 13632
rect 11614 13572 11618 13628
rect 11618 13572 11674 13628
rect 11674 13572 11678 13628
rect 11614 13568 11678 13572
rect 18322 13628 18386 13632
rect 18322 13572 18326 13628
rect 18326 13572 18382 13628
rect 18382 13572 18386 13628
rect 18322 13568 18386 13572
rect 18402 13628 18466 13632
rect 18402 13572 18406 13628
rect 18406 13572 18462 13628
rect 18462 13572 18466 13628
rect 18402 13568 18466 13572
rect 18482 13628 18546 13632
rect 18482 13572 18486 13628
rect 18486 13572 18542 13628
rect 18542 13572 18546 13628
rect 18482 13568 18546 13572
rect 18562 13628 18626 13632
rect 18562 13572 18566 13628
rect 18566 13572 18622 13628
rect 18622 13572 18626 13628
rect 18562 13568 18626 13572
rect 25270 13628 25334 13632
rect 25270 13572 25274 13628
rect 25274 13572 25330 13628
rect 25330 13572 25334 13628
rect 25270 13568 25334 13572
rect 25350 13628 25414 13632
rect 25350 13572 25354 13628
rect 25354 13572 25410 13628
rect 25410 13572 25414 13628
rect 25350 13568 25414 13572
rect 25430 13628 25494 13632
rect 25430 13572 25434 13628
rect 25434 13572 25490 13628
rect 25490 13572 25494 13628
rect 25430 13568 25494 13572
rect 25510 13628 25574 13632
rect 25510 13572 25514 13628
rect 25514 13572 25570 13628
rect 25570 13572 25574 13628
rect 25510 13568 25574 13572
rect 7900 13084 7964 13088
rect 7900 13028 7904 13084
rect 7904 13028 7960 13084
rect 7960 13028 7964 13084
rect 7900 13024 7964 13028
rect 7980 13084 8044 13088
rect 7980 13028 7984 13084
rect 7984 13028 8040 13084
rect 8040 13028 8044 13084
rect 7980 13024 8044 13028
rect 8060 13084 8124 13088
rect 8060 13028 8064 13084
rect 8064 13028 8120 13084
rect 8120 13028 8124 13084
rect 8060 13024 8124 13028
rect 8140 13084 8204 13088
rect 8140 13028 8144 13084
rect 8144 13028 8200 13084
rect 8200 13028 8204 13084
rect 8140 13024 8204 13028
rect 14848 13084 14912 13088
rect 14848 13028 14852 13084
rect 14852 13028 14908 13084
rect 14908 13028 14912 13084
rect 14848 13024 14912 13028
rect 14928 13084 14992 13088
rect 14928 13028 14932 13084
rect 14932 13028 14988 13084
rect 14988 13028 14992 13084
rect 14928 13024 14992 13028
rect 15008 13084 15072 13088
rect 15008 13028 15012 13084
rect 15012 13028 15068 13084
rect 15068 13028 15072 13084
rect 15008 13024 15072 13028
rect 15088 13084 15152 13088
rect 15088 13028 15092 13084
rect 15092 13028 15148 13084
rect 15148 13028 15152 13084
rect 15088 13024 15152 13028
rect 21796 13084 21860 13088
rect 21796 13028 21800 13084
rect 21800 13028 21856 13084
rect 21856 13028 21860 13084
rect 21796 13024 21860 13028
rect 21876 13084 21940 13088
rect 21876 13028 21880 13084
rect 21880 13028 21936 13084
rect 21936 13028 21940 13084
rect 21876 13024 21940 13028
rect 21956 13084 22020 13088
rect 21956 13028 21960 13084
rect 21960 13028 22016 13084
rect 22016 13028 22020 13084
rect 21956 13024 22020 13028
rect 22036 13084 22100 13088
rect 22036 13028 22040 13084
rect 22040 13028 22096 13084
rect 22096 13028 22100 13084
rect 22036 13024 22100 13028
rect 4426 12540 4490 12544
rect 4426 12484 4430 12540
rect 4430 12484 4486 12540
rect 4486 12484 4490 12540
rect 4426 12480 4490 12484
rect 4506 12540 4570 12544
rect 4506 12484 4510 12540
rect 4510 12484 4566 12540
rect 4566 12484 4570 12540
rect 4506 12480 4570 12484
rect 4586 12540 4650 12544
rect 4586 12484 4590 12540
rect 4590 12484 4646 12540
rect 4646 12484 4650 12540
rect 4586 12480 4650 12484
rect 4666 12540 4730 12544
rect 4666 12484 4670 12540
rect 4670 12484 4726 12540
rect 4726 12484 4730 12540
rect 4666 12480 4730 12484
rect 11374 12540 11438 12544
rect 11374 12484 11378 12540
rect 11378 12484 11434 12540
rect 11434 12484 11438 12540
rect 11374 12480 11438 12484
rect 11454 12540 11518 12544
rect 11454 12484 11458 12540
rect 11458 12484 11514 12540
rect 11514 12484 11518 12540
rect 11454 12480 11518 12484
rect 11534 12540 11598 12544
rect 11534 12484 11538 12540
rect 11538 12484 11594 12540
rect 11594 12484 11598 12540
rect 11534 12480 11598 12484
rect 11614 12540 11678 12544
rect 11614 12484 11618 12540
rect 11618 12484 11674 12540
rect 11674 12484 11678 12540
rect 11614 12480 11678 12484
rect 18322 12540 18386 12544
rect 18322 12484 18326 12540
rect 18326 12484 18382 12540
rect 18382 12484 18386 12540
rect 18322 12480 18386 12484
rect 18402 12540 18466 12544
rect 18402 12484 18406 12540
rect 18406 12484 18462 12540
rect 18462 12484 18466 12540
rect 18402 12480 18466 12484
rect 18482 12540 18546 12544
rect 18482 12484 18486 12540
rect 18486 12484 18542 12540
rect 18542 12484 18546 12540
rect 18482 12480 18546 12484
rect 18562 12540 18626 12544
rect 18562 12484 18566 12540
rect 18566 12484 18622 12540
rect 18622 12484 18626 12540
rect 18562 12480 18626 12484
rect 25270 12540 25334 12544
rect 25270 12484 25274 12540
rect 25274 12484 25330 12540
rect 25330 12484 25334 12540
rect 25270 12480 25334 12484
rect 25350 12540 25414 12544
rect 25350 12484 25354 12540
rect 25354 12484 25410 12540
rect 25410 12484 25414 12540
rect 25350 12480 25414 12484
rect 25430 12540 25494 12544
rect 25430 12484 25434 12540
rect 25434 12484 25490 12540
rect 25490 12484 25494 12540
rect 25430 12480 25494 12484
rect 25510 12540 25574 12544
rect 25510 12484 25514 12540
rect 25514 12484 25570 12540
rect 25570 12484 25574 12540
rect 25510 12480 25574 12484
rect 7900 11996 7964 12000
rect 7900 11940 7904 11996
rect 7904 11940 7960 11996
rect 7960 11940 7964 11996
rect 7900 11936 7964 11940
rect 7980 11996 8044 12000
rect 7980 11940 7984 11996
rect 7984 11940 8040 11996
rect 8040 11940 8044 11996
rect 7980 11936 8044 11940
rect 8060 11996 8124 12000
rect 8060 11940 8064 11996
rect 8064 11940 8120 11996
rect 8120 11940 8124 11996
rect 8060 11936 8124 11940
rect 8140 11996 8204 12000
rect 8140 11940 8144 11996
rect 8144 11940 8200 11996
rect 8200 11940 8204 11996
rect 8140 11936 8204 11940
rect 14848 11996 14912 12000
rect 14848 11940 14852 11996
rect 14852 11940 14908 11996
rect 14908 11940 14912 11996
rect 14848 11936 14912 11940
rect 14928 11996 14992 12000
rect 14928 11940 14932 11996
rect 14932 11940 14988 11996
rect 14988 11940 14992 11996
rect 14928 11936 14992 11940
rect 15008 11996 15072 12000
rect 15008 11940 15012 11996
rect 15012 11940 15068 11996
rect 15068 11940 15072 11996
rect 15008 11936 15072 11940
rect 15088 11996 15152 12000
rect 15088 11940 15092 11996
rect 15092 11940 15148 11996
rect 15148 11940 15152 11996
rect 15088 11936 15152 11940
rect 21796 11996 21860 12000
rect 21796 11940 21800 11996
rect 21800 11940 21856 11996
rect 21856 11940 21860 11996
rect 21796 11936 21860 11940
rect 21876 11996 21940 12000
rect 21876 11940 21880 11996
rect 21880 11940 21936 11996
rect 21936 11940 21940 11996
rect 21876 11936 21940 11940
rect 21956 11996 22020 12000
rect 21956 11940 21960 11996
rect 21960 11940 22016 11996
rect 22016 11940 22020 11996
rect 21956 11936 22020 11940
rect 22036 11996 22100 12000
rect 22036 11940 22040 11996
rect 22040 11940 22096 11996
rect 22096 11940 22100 11996
rect 22036 11936 22100 11940
rect 4426 11452 4490 11456
rect 4426 11396 4430 11452
rect 4430 11396 4486 11452
rect 4486 11396 4490 11452
rect 4426 11392 4490 11396
rect 4506 11452 4570 11456
rect 4506 11396 4510 11452
rect 4510 11396 4566 11452
rect 4566 11396 4570 11452
rect 4506 11392 4570 11396
rect 4586 11452 4650 11456
rect 4586 11396 4590 11452
rect 4590 11396 4646 11452
rect 4646 11396 4650 11452
rect 4586 11392 4650 11396
rect 4666 11452 4730 11456
rect 4666 11396 4670 11452
rect 4670 11396 4726 11452
rect 4726 11396 4730 11452
rect 4666 11392 4730 11396
rect 11374 11452 11438 11456
rect 11374 11396 11378 11452
rect 11378 11396 11434 11452
rect 11434 11396 11438 11452
rect 11374 11392 11438 11396
rect 11454 11452 11518 11456
rect 11454 11396 11458 11452
rect 11458 11396 11514 11452
rect 11514 11396 11518 11452
rect 11454 11392 11518 11396
rect 11534 11452 11598 11456
rect 11534 11396 11538 11452
rect 11538 11396 11594 11452
rect 11594 11396 11598 11452
rect 11534 11392 11598 11396
rect 11614 11452 11678 11456
rect 11614 11396 11618 11452
rect 11618 11396 11674 11452
rect 11674 11396 11678 11452
rect 11614 11392 11678 11396
rect 18322 11452 18386 11456
rect 18322 11396 18326 11452
rect 18326 11396 18382 11452
rect 18382 11396 18386 11452
rect 18322 11392 18386 11396
rect 18402 11452 18466 11456
rect 18402 11396 18406 11452
rect 18406 11396 18462 11452
rect 18462 11396 18466 11452
rect 18402 11392 18466 11396
rect 18482 11452 18546 11456
rect 18482 11396 18486 11452
rect 18486 11396 18542 11452
rect 18542 11396 18546 11452
rect 18482 11392 18546 11396
rect 18562 11452 18626 11456
rect 18562 11396 18566 11452
rect 18566 11396 18622 11452
rect 18622 11396 18626 11452
rect 18562 11392 18626 11396
rect 25270 11452 25334 11456
rect 25270 11396 25274 11452
rect 25274 11396 25330 11452
rect 25330 11396 25334 11452
rect 25270 11392 25334 11396
rect 25350 11452 25414 11456
rect 25350 11396 25354 11452
rect 25354 11396 25410 11452
rect 25410 11396 25414 11452
rect 25350 11392 25414 11396
rect 25430 11452 25494 11456
rect 25430 11396 25434 11452
rect 25434 11396 25490 11452
rect 25490 11396 25494 11452
rect 25430 11392 25494 11396
rect 25510 11452 25574 11456
rect 25510 11396 25514 11452
rect 25514 11396 25570 11452
rect 25570 11396 25574 11452
rect 25510 11392 25574 11396
rect 7900 10908 7964 10912
rect 7900 10852 7904 10908
rect 7904 10852 7960 10908
rect 7960 10852 7964 10908
rect 7900 10848 7964 10852
rect 7980 10908 8044 10912
rect 7980 10852 7984 10908
rect 7984 10852 8040 10908
rect 8040 10852 8044 10908
rect 7980 10848 8044 10852
rect 8060 10908 8124 10912
rect 8060 10852 8064 10908
rect 8064 10852 8120 10908
rect 8120 10852 8124 10908
rect 8060 10848 8124 10852
rect 8140 10908 8204 10912
rect 8140 10852 8144 10908
rect 8144 10852 8200 10908
rect 8200 10852 8204 10908
rect 8140 10848 8204 10852
rect 14848 10908 14912 10912
rect 14848 10852 14852 10908
rect 14852 10852 14908 10908
rect 14908 10852 14912 10908
rect 14848 10848 14912 10852
rect 14928 10908 14992 10912
rect 14928 10852 14932 10908
rect 14932 10852 14988 10908
rect 14988 10852 14992 10908
rect 14928 10848 14992 10852
rect 15008 10908 15072 10912
rect 15008 10852 15012 10908
rect 15012 10852 15068 10908
rect 15068 10852 15072 10908
rect 15008 10848 15072 10852
rect 15088 10908 15152 10912
rect 15088 10852 15092 10908
rect 15092 10852 15148 10908
rect 15148 10852 15152 10908
rect 15088 10848 15152 10852
rect 21796 10908 21860 10912
rect 21796 10852 21800 10908
rect 21800 10852 21856 10908
rect 21856 10852 21860 10908
rect 21796 10848 21860 10852
rect 21876 10908 21940 10912
rect 21876 10852 21880 10908
rect 21880 10852 21936 10908
rect 21936 10852 21940 10908
rect 21876 10848 21940 10852
rect 21956 10908 22020 10912
rect 21956 10852 21960 10908
rect 21960 10852 22016 10908
rect 22016 10852 22020 10908
rect 21956 10848 22020 10852
rect 22036 10908 22100 10912
rect 22036 10852 22040 10908
rect 22040 10852 22096 10908
rect 22096 10852 22100 10908
rect 22036 10848 22100 10852
rect 4426 10364 4490 10368
rect 4426 10308 4430 10364
rect 4430 10308 4486 10364
rect 4486 10308 4490 10364
rect 4426 10304 4490 10308
rect 4506 10364 4570 10368
rect 4506 10308 4510 10364
rect 4510 10308 4566 10364
rect 4566 10308 4570 10364
rect 4506 10304 4570 10308
rect 4586 10364 4650 10368
rect 4586 10308 4590 10364
rect 4590 10308 4646 10364
rect 4646 10308 4650 10364
rect 4586 10304 4650 10308
rect 4666 10364 4730 10368
rect 4666 10308 4670 10364
rect 4670 10308 4726 10364
rect 4726 10308 4730 10364
rect 4666 10304 4730 10308
rect 11374 10364 11438 10368
rect 11374 10308 11378 10364
rect 11378 10308 11434 10364
rect 11434 10308 11438 10364
rect 11374 10304 11438 10308
rect 11454 10364 11518 10368
rect 11454 10308 11458 10364
rect 11458 10308 11514 10364
rect 11514 10308 11518 10364
rect 11454 10304 11518 10308
rect 11534 10364 11598 10368
rect 11534 10308 11538 10364
rect 11538 10308 11594 10364
rect 11594 10308 11598 10364
rect 11534 10304 11598 10308
rect 11614 10364 11678 10368
rect 11614 10308 11618 10364
rect 11618 10308 11674 10364
rect 11674 10308 11678 10364
rect 11614 10304 11678 10308
rect 18322 10364 18386 10368
rect 18322 10308 18326 10364
rect 18326 10308 18382 10364
rect 18382 10308 18386 10364
rect 18322 10304 18386 10308
rect 18402 10364 18466 10368
rect 18402 10308 18406 10364
rect 18406 10308 18462 10364
rect 18462 10308 18466 10364
rect 18402 10304 18466 10308
rect 18482 10364 18546 10368
rect 18482 10308 18486 10364
rect 18486 10308 18542 10364
rect 18542 10308 18546 10364
rect 18482 10304 18546 10308
rect 18562 10364 18626 10368
rect 18562 10308 18566 10364
rect 18566 10308 18622 10364
rect 18622 10308 18626 10364
rect 18562 10304 18626 10308
rect 25270 10364 25334 10368
rect 25270 10308 25274 10364
rect 25274 10308 25330 10364
rect 25330 10308 25334 10364
rect 25270 10304 25334 10308
rect 25350 10364 25414 10368
rect 25350 10308 25354 10364
rect 25354 10308 25410 10364
rect 25410 10308 25414 10364
rect 25350 10304 25414 10308
rect 25430 10364 25494 10368
rect 25430 10308 25434 10364
rect 25434 10308 25490 10364
rect 25490 10308 25494 10364
rect 25430 10304 25494 10308
rect 25510 10364 25574 10368
rect 25510 10308 25514 10364
rect 25514 10308 25570 10364
rect 25570 10308 25574 10364
rect 25510 10304 25574 10308
rect 7900 9820 7964 9824
rect 7900 9764 7904 9820
rect 7904 9764 7960 9820
rect 7960 9764 7964 9820
rect 7900 9760 7964 9764
rect 7980 9820 8044 9824
rect 7980 9764 7984 9820
rect 7984 9764 8040 9820
rect 8040 9764 8044 9820
rect 7980 9760 8044 9764
rect 8060 9820 8124 9824
rect 8060 9764 8064 9820
rect 8064 9764 8120 9820
rect 8120 9764 8124 9820
rect 8060 9760 8124 9764
rect 8140 9820 8204 9824
rect 8140 9764 8144 9820
rect 8144 9764 8200 9820
rect 8200 9764 8204 9820
rect 8140 9760 8204 9764
rect 14848 9820 14912 9824
rect 14848 9764 14852 9820
rect 14852 9764 14908 9820
rect 14908 9764 14912 9820
rect 14848 9760 14912 9764
rect 14928 9820 14992 9824
rect 14928 9764 14932 9820
rect 14932 9764 14988 9820
rect 14988 9764 14992 9820
rect 14928 9760 14992 9764
rect 15008 9820 15072 9824
rect 15008 9764 15012 9820
rect 15012 9764 15068 9820
rect 15068 9764 15072 9820
rect 15008 9760 15072 9764
rect 15088 9820 15152 9824
rect 15088 9764 15092 9820
rect 15092 9764 15148 9820
rect 15148 9764 15152 9820
rect 15088 9760 15152 9764
rect 21796 9820 21860 9824
rect 21796 9764 21800 9820
rect 21800 9764 21856 9820
rect 21856 9764 21860 9820
rect 21796 9760 21860 9764
rect 21876 9820 21940 9824
rect 21876 9764 21880 9820
rect 21880 9764 21936 9820
rect 21936 9764 21940 9820
rect 21876 9760 21940 9764
rect 21956 9820 22020 9824
rect 21956 9764 21960 9820
rect 21960 9764 22016 9820
rect 22016 9764 22020 9820
rect 21956 9760 22020 9764
rect 22036 9820 22100 9824
rect 22036 9764 22040 9820
rect 22040 9764 22096 9820
rect 22096 9764 22100 9820
rect 22036 9760 22100 9764
rect 4426 9276 4490 9280
rect 4426 9220 4430 9276
rect 4430 9220 4486 9276
rect 4486 9220 4490 9276
rect 4426 9216 4490 9220
rect 4506 9276 4570 9280
rect 4506 9220 4510 9276
rect 4510 9220 4566 9276
rect 4566 9220 4570 9276
rect 4506 9216 4570 9220
rect 4586 9276 4650 9280
rect 4586 9220 4590 9276
rect 4590 9220 4646 9276
rect 4646 9220 4650 9276
rect 4586 9216 4650 9220
rect 4666 9276 4730 9280
rect 4666 9220 4670 9276
rect 4670 9220 4726 9276
rect 4726 9220 4730 9276
rect 4666 9216 4730 9220
rect 11374 9276 11438 9280
rect 11374 9220 11378 9276
rect 11378 9220 11434 9276
rect 11434 9220 11438 9276
rect 11374 9216 11438 9220
rect 11454 9276 11518 9280
rect 11454 9220 11458 9276
rect 11458 9220 11514 9276
rect 11514 9220 11518 9276
rect 11454 9216 11518 9220
rect 11534 9276 11598 9280
rect 11534 9220 11538 9276
rect 11538 9220 11594 9276
rect 11594 9220 11598 9276
rect 11534 9216 11598 9220
rect 11614 9276 11678 9280
rect 11614 9220 11618 9276
rect 11618 9220 11674 9276
rect 11674 9220 11678 9276
rect 11614 9216 11678 9220
rect 18322 9276 18386 9280
rect 18322 9220 18326 9276
rect 18326 9220 18382 9276
rect 18382 9220 18386 9276
rect 18322 9216 18386 9220
rect 18402 9276 18466 9280
rect 18402 9220 18406 9276
rect 18406 9220 18462 9276
rect 18462 9220 18466 9276
rect 18402 9216 18466 9220
rect 18482 9276 18546 9280
rect 18482 9220 18486 9276
rect 18486 9220 18542 9276
rect 18542 9220 18546 9276
rect 18482 9216 18546 9220
rect 18562 9276 18626 9280
rect 18562 9220 18566 9276
rect 18566 9220 18622 9276
rect 18622 9220 18626 9276
rect 18562 9216 18626 9220
rect 25270 9276 25334 9280
rect 25270 9220 25274 9276
rect 25274 9220 25330 9276
rect 25330 9220 25334 9276
rect 25270 9216 25334 9220
rect 25350 9276 25414 9280
rect 25350 9220 25354 9276
rect 25354 9220 25410 9276
rect 25410 9220 25414 9276
rect 25350 9216 25414 9220
rect 25430 9276 25494 9280
rect 25430 9220 25434 9276
rect 25434 9220 25490 9276
rect 25490 9220 25494 9276
rect 25430 9216 25494 9220
rect 25510 9276 25574 9280
rect 25510 9220 25514 9276
rect 25514 9220 25570 9276
rect 25570 9220 25574 9276
rect 25510 9216 25574 9220
rect 7900 8732 7964 8736
rect 7900 8676 7904 8732
rect 7904 8676 7960 8732
rect 7960 8676 7964 8732
rect 7900 8672 7964 8676
rect 7980 8732 8044 8736
rect 7980 8676 7984 8732
rect 7984 8676 8040 8732
rect 8040 8676 8044 8732
rect 7980 8672 8044 8676
rect 8060 8732 8124 8736
rect 8060 8676 8064 8732
rect 8064 8676 8120 8732
rect 8120 8676 8124 8732
rect 8060 8672 8124 8676
rect 8140 8732 8204 8736
rect 8140 8676 8144 8732
rect 8144 8676 8200 8732
rect 8200 8676 8204 8732
rect 8140 8672 8204 8676
rect 14848 8732 14912 8736
rect 14848 8676 14852 8732
rect 14852 8676 14908 8732
rect 14908 8676 14912 8732
rect 14848 8672 14912 8676
rect 14928 8732 14992 8736
rect 14928 8676 14932 8732
rect 14932 8676 14988 8732
rect 14988 8676 14992 8732
rect 14928 8672 14992 8676
rect 15008 8732 15072 8736
rect 15008 8676 15012 8732
rect 15012 8676 15068 8732
rect 15068 8676 15072 8732
rect 15008 8672 15072 8676
rect 15088 8732 15152 8736
rect 15088 8676 15092 8732
rect 15092 8676 15148 8732
rect 15148 8676 15152 8732
rect 15088 8672 15152 8676
rect 21796 8732 21860 8736
rect 21796 8676 21800 8732
rect 21800 8676 21856 8732
rect 21856 8676 21860 8732
rect 21796 8672 21860 8676
rect 21876 8732 21940 8736
rect 21876 8676 21880 8732
rect 21880 8676 21936 8732
rect 21936 8676 21940 8732
rect 21876 8672 21940 8676
rect 21956 8732 22020 8736
rect 21956 8676 21960 8732
rect 21960 8676 22016 8732
rect 22016 8676 22020 8732
rect 21956 8672 22020 8676
rect 22036 8732 22100 8736
rect 22036 8676 22040 8732
rect 22040 8676 22096 8732
rect 22096 8676 22100 8732
rect 22036 8672 22100 8676
rect 4426 8188 4490 8192
rect 4426 8132 4430 8188
rect 4430 8132 4486 8188
rect 4486 8132 4490 8188
rect 4426 8128 4490 8132
rect 4506 8188 4570 8192
rect 4506 8132 4510 8188
rect 4510 8132 4566 8188
rect 4566 8132 4570 8188
rect 4506 8128 4570 8132
rect 4586 8188 4650 8192
rect 4586 8132 4590 8188
rect 4590 8132 4646 8188
rect 4646 8132 4650 8188
rect 4586 8128 4650 8132
rect 4666 8188 4730 8192
rect 4666 8132 4670 8188
rect 4670 8132 4726 8188
rect 4726 8132 4730 8188
rect 4666 8128 4730 8132
rect 11374 8188 11438 8192
rect 11374 8132 11378 8188
rect 11378 8132 11434 8188
rect 11434 8132 11438 8188
rect 11374 8128 11438 8132
rect 11454 8188 11518 8192
rect 11454 8132 11458 8188
rect 11458 8132 11514 8188
rect 11514 8132 11518 8188
rect 11454 8128 11518 8132
rect 11534 8188 11598 8192
rect 11534 8132 11538 8188
rect 11538 8132 11594 8188
rect 11594 8132 11598 8188
rect 11534 8128 11598 8132
rect 11614 8188 11678 8192
rect 11614 8132 11618 8188
rect 11618 8132 11674 8188
rect 11674 8132 11678 8188
rect 11614 8128 11678 8132
rect 18322 8188 18386 8192
rect 18322 8132 18326 8188
rect 18326 8132 18382 8188
rect 18382 8132 18386 8188
rect 18322 8128 18386 8132
rect 18402 8188 18466 8192
rect 18402 8132 18406 8188
rect 18406 8132 18462 8188
rect 18462 8132 18466 8188
rect 18402 8128 18466 8132
rect 18482 8188 18546 8192
rect 18482 8132 18486 8188
rect 18486 8132 18542 8188
rect 18542 8132 18546 8188
rect 18482 8128 18546 8132
rect 18562 8188 18626 8192
rect 18562 8132 18566 8188
rect 18566 8132 18622 8188
rect 18622 8132 18626 8188
rect 18562 8128 18626 8132
rect 25270 8188 25334 8192
rect 25270 8132 25274 8188
rect 25274 8132 25330 8188
rect 25330 8132 25334 8188
rect 25270 8128 25334 8132
rect 25350 8188 25414 8192
rect 25350 8132 25354 8188
rect 25354 8132 25410 8188
rect 25410 8132 25414 8188
rect 25350 8128 25414 8132
rect 25430 8188 25494 8192
rect 25430 8132 25434 8188
rect 25434 8132 25490 8188
rect 25490 8132 25494 8188
rect 25430 8128 25494 8132
rect 25510 8188 25574 8192
rect 25510 8132 25514 8188
rect 25514 8132 25570 8188
rect 25570 8132 25574 8188
rect 25510 8128 25574 8132
rect 7900 7644 7964 7648
rect 7900 7588 7904 7644
rect 7904 7588 7960 7644
rect 7960 7588 7964 7644
rect 7900 7584 7964 7588
rect 7980 7644 8044 7648
rect 7980 7588 7984 7644
rect 7984 7588 8040 7644
rect 8040 7588 8044 7644
rect 7980 7584 8044 7588
rect 8060 7644 8124 7648
rect 8060 7588 8064 7644
rect 8064 7588 8120 7644
rect 8120 7588 8124 7644
rect 8060 7584 8124 7588
rect 8140 7644 8204 7648
rect 8140 7588 8144 7644
rect 8144 7588 8200 7644
rect 8200 7588 8204 7644
rect 8140 7584 8204 7588
rect 14848 7644 14912 7648
rect 14848 7588 14852 7644
rect 14852 7588 14908 7644
rect 14908 7588 14912 7644
rect 14848 7584 14912 7588
rect 14928 7644 14992 7648
rect 14928 7588 14932 7644
rect 14932 7588 14988 7644
rect 14988 7588 14992 7644
rect 14928 7584 14992 7588
rect 15008 7644 15072 7648
rect 15008 7588 15012 7644
rect 15012 7588 15068 7644
rect 15068 7588 15072 7644
rect 15008 7584 15072 7588
rect 15088 7644 15152 7648
rect 15088 7588 15092 7644
rect 15092 7588 15148 7644
rect 15148 7588 15152 7644
rect 15088 7584 15152 7588
rect 21796 7644 21860 7648
rect 21796 7588 21800 7644
rect 21800 7588 21856 7644
rect 21856 7588 21860 7644
rect 21796 7584 21860 7588
rect 21876 7644 21940 7648
rect 21876 7588 21880 7644
rect 21880 7588 21936 7644
rect 21936 7588 21940 7644
rect 21876 7584 21940 7588
rect 21956 7644 22020 7648
rect 21956 7588 21960 7644
rect 21960 7588 22016 7644
rect 22016 7588 22020 7644
rect 21956 7584 22020 7588
rect 22036 7644 22100 7648
rect 22036 7588 22040 7644
rect 22040 7588 22096 7644
rect 22096 7588 22100 7644
rect 22036 7584 22100 7588
rect 4426 7100 4490 7104
rect 4426 7044 4430 7100
rect 4430 7044 4486 7100
rect 4486 7044 4490 7100
rect 4426 7040 4490 7044
rect 4506 7100 4570 7104
rect 4506 7044 4510 7100
rect 4510 7044 4566 7100
rect 4566 7044 4570 7100
rect 4506 7040 4570 7044
rect 4586 7100 4650 7104
rect 4586 7044 4590 7100
rect 4590 7044 4646 7100
rect 4646 7044 4650 7100
rect 4586 7040 4650 7044
rect 4666 7100 4730 7104
rect 4666 7044 4670 7100
rect 4670 7044 4726 7100
rect 4726 7044 4730 7100
rect 4666 7040 4730 7044
rect 11374 7100 11438 7104
rect 11374 7044 11378 7100
rect 11378 7044 11434 7100
rect 11434 7044 11438 7100
rect 11374 7040 11438 7044
rect 11454 7100 11518 7104
rect 11454 7044 11458 7100
rect 11458 7044 11514 7100
rect 11514 7044 11518 7100
rect 11454 7040 11518 7044
rect 11534 7100 11598 7104
rect 11534 7044 11538 7100
rect 11538 7044 11594 7100
rect 11594 7044 11598 7100
rect 11534 7040 11598 7044
rect 11614 7100 11678 7104
rect 11614 7044 11618 7100
rect 11618 7044 11674 7100
rect 11674 7044 11678 7100
rect 11614 7040 11678 7044
rect 18322 7100 18386 7104
rect 18322 7044 18326 7100
rect 18326 7044 18382 7100
rect 18382 7044 18386 7100
rect 18322 7040 18386 7044
rect 18402 7100 18466 7104
rect 18402 7044 18406 7100
rect 18406 7044 18462 7100
rect 18462 7044 18466 7100
rect 18402 7040 18466 7044
rect 18482 7100 18546 7104
rect 18482 7044 18486 7100
rect 18486 7044 18542 7100
rect 18542 7044 18546 7100
rect 18482 7040 18546 7044
rect 18562 7100 18626 7104
rect 18562 7044 18566 7100
rect 18566 7044 18622 7100
rect 18622 7044 18626 7100
rect 18562 7040 18626 7044
rect 25270 7100 25334 7104
rect 25270 7044 25274 7100
rect 25274 7044 25330 7100
rect 25330 7044 25334 7100
rect 25270 7040 25334 7044
rect 25350 7100 25414 7104
rect 25350 7044 25354 7100
rect 25354 7044 25410 7100
rect 25410 7044 25414 7100
rect 25350 7040 25414 7044
rect 25430 7100 25494 7104
rect 25430 7044 25434 7100
rect 25434 7044 25490 7100
rect 25490 7044 25494 7100
rect 25430 7040 25494 7044
rect 25510 7100 25574 7104
rect 25510 7044 25514 7100
rect 25514 7044 25570 7100
rect 25570 7044 25574 7100
rect 25510 7040 25574 7044
rect 7900 6556 7964 6560
rect 7900 6500 7904 6556
rect 7904 6500 7960 6556
rect 7960 6500 7964 6556
rect 7900 6496 7964 6500
rect 7980 6556 8044 6560
rect 7980 6500 7984 6556
rect 7984 6500 8040 6556
rect 8040 6500 8044 6556
rect 7980 6496 8044 6500
rect 8060 6556 8124 6560
rect 8060 6500 8064 6556
rect 8064 6500 8120 6556
rect 8120 6500 8124 6556
rect 8060 6496 8124 6500
rect 8140 6556 8204 6560
rect 8140 6500 8144 6556
rect 8144 6500 8200 6556
rect 8200 6500 8204 6556
rect 8140 6496 8204 6500
rect 14848 6556 14912 6560
rect 14848 6500 14852 6556
rect 14852 6500 14908 6556
rect 14908 6500 14912 6556
rect 14848 6496 14912 6500
rect 14928 6556 14992 6560
rect 14928 6500 14932 6556
rect 14932 6500 14988 6556
rect 14988 6500 14992 6556
rect 14928 6496 14992 6500
rect 15008 6556 15072 6560
rect 15008 6500 15012 6556
rect 15012 6500 15068 6556
rect 15068 6500 15072 6556
rect 15008 6496 15072 6500
rect 15088 6556 15152 6560
rect 15088 6500 15092 6556
rect 15092 6500 15148 6556
rect 15148 6500 15152 6556
rect 15088 6496 15152 6500
rect 21796 6556 21860 6560
rect 21796 6500 21800 6556
rect 21800 6500 21856 6556
rect 21856 6500 21860 6556
rect 21796 6496 21860 6500
rect 21876 6556 21940 6560
rect 21876 6500 21880 6556
rect 21880 6500 21936 6556
rect 21936 6500 21940 6556
rect 21876 6496 21940 6500
rect 21956 6556 22020 6560
rect 21956 6500 21960 6556
rect 21960 6500 22016 6556
rect 22016 6500 22020 6556
rect 21956 6496 22020 6500
rect 22036 6556 22100 6560
rect 22036 6500 22040 6556
rect 22040 6500 22096 6556
rect 22096 6500 22100 6556
rect 22036 6496 22100 6500
rect 4426 6012 4490 6016
rect 4426 5956 4430 6012
rect 4430 5956 4486 6012
rect 4486 5956 4490 6012
rect 4426 5952 4490 5956
rect 4506 6012 4570 6016
rect 4506 5956 4510 6012
rect 4510 5956 4566 6012
rect 4566 5956 4570 6012
rect 4506 5952 4570 5956
rect 4586 6012 4650 6016
rect 4586 5956 4590 6012
rect 4590 5956 4646 6012
rect 4646 5956 4650 6012
rect 4586 5952 4650 5956
rect 4666 6012 4730 6016
rect 4666 5956 4670 6012
rect 4670 5956 4726 6012
rect 4726 5956 4730 6012
rect 4666 5952 4730 5956
rect 11374 6012 11438 6016
rect 11374 5956 11378 6012
rect 11378 5956 11434 6012
rect 11434 5956 11438 6012
rect 11374 5952 11438 5956
rect 11454 6012 11518 6016
rect 11454 5956 11458 6012
rect 11458 5956 11514 6012
rect 11514 5956 11518 6012
rect 11454 5952 11518 5956
rect 11534 6012 11598 6016
rect 11534 5956 11538 6012
rect 11538 5956 11594 6012
rect 11594 5956 11598 6012
rect 11534 5952 11598 5956
rect 11614 6012 11678 6016
rect 11614 5956 11618 6012
rect 11618 5956 11674 6012
rect 11674 5956 11678 6012
rect 11614 5952 11678 5956
rect 18322 6012 18386 6016
rect 18322 5956 18326 6012
rect 18326 5956 18382 6012
rect 18382 5956 18386 6012
rect 18322 5952 18386 5956
rect 18402 6012 18466 6016
rect 18402 5956 18406 6012
rect 18406 5956 18462 6012
rect 18462 5956 18466 6012
rect 18402 5952 18466 5956
rect 18482 6012 18546 6016
rect 18482 5956 18486 6012
rect 18486 5956 18542 6012
rect 18542 5956 18546 6012
rect 18482 5952 18546 5956
rect 18562 6012 18626 6016
rect 18562 5956 18566 6012
rect 18566 5956 18622 6012
rect 18622 5956 18626 6012
rect 18562 5952 18626 5956
rect 25270 6012 25334 6016
rect 25270 5956 25274 6012
rect 25274 5956 25330 6012
rect 25330 5956 25334 6012
rect 25270 5952 25334 5956
rect 25350 6012 25414 6016
rect 25350 5956 25354 6012
rect 25354 5956 25410 6012
rect 25410 5956 25414 6012
rect 25350 5952 25414 5956
rect 25430 6012 25494 6016
rect 25430 5956 25434 6012
rect 25434 5956 25490 6012
rect 25490 5956 25494 6012
rect 25430 5952 25494 5956
rect 25510 6012 25574 6016
rect 25510 5956 25514 6012
rect 25514 5956 25570 6012
rect 25570 5956 25574 6012
rect 25510 5952 25574 5956
rect 7900 5468 7964 5472
rect 7900 5412 7904 5468
rect 7904 5412 7960 5468
rect 7960 5412 7964 5468
rect 7900 5408 7964 5412
rect 7980 5468 8044 5472
rect 7980 5412 7984 5468
rect 7984 5412 8040 5468
rect 8040 5412 8044 5468
rect 7980 5408 8044 5412
rect 8060 5468 8124 5472
rect 8060 5412 8064 5468
rect 8064 5412 8120 5468
rect 8120 5412 8124 5468
rect 8060 5408 8124 5412
rect 8140 5468 8204 5472
rect 8140 5412 8144 5468
rect 8144 5412 8200 5468
rect 8200 5412 8204 5468
rect 8140 5408 8204 5412
rect 14848 5468 14912 5472
rect 14848 5412 14852 5468
rect 14852 5412 14908 5468
rect 14908 5412 14912 5468
rect 14848 5408 14912 5412
rect 14928 5468 14992 5472
rect 14928 5412 14932 5468
rect 14932 5412 14988 5468
rect 14988 5412 14992 5468
rect 14928 5408 14992 5412
rect 15008 5468 15072 5472
rect 15008 5412 15012 5468
rect 15012 5412 15068 5468
rect 15068 5412 15072 5468
rect 15008 5408 15072 5412
rect 15088 5468 15152 5472
rect 15088 5412 15092 5468
rect 15092 5412 15148 5468
rect 15148 5412 15152 5468
rect 15088 5408 15152 5412
rect 21796 5468 21860 5472
rect 21796 5412 21800 5468
rect 21800 5412 21856 5468
rect 21856 5412 21860 5468
rect 21796 5408 21860 5412
rect 21876 5468 21940 5472
rect 21876 5412 21880 5468
rect 21880 5412 21936 5468
rect 21936 5412 21940 5468
rect 21876 5408 21940 5412
rect 21956 5468 22020 5472
rect 21956 5412 21960 5468
rect 21960 5412 22016 5468
rect 22016 5412 22020 5468
rect 21956 5408 22020 5412
rect 22036 5468 22100 5472
rect 22036 5412 22040 5468
rect 22040 5412 22096 5468
rect 22096 5412 22100 5468
rect 22036 5408 22100 5412
rect 4426 4924 4490 4928
rect 4426 4868 4430 4924
rect 4430 4868 4486 4924
rect 4486 4868 4490 4924
rect 4426 4864 4490 4868
rect 4506 4924 4570 4928
rect 4506 4868 4510 4924
rect 4510 4868 4566 4924
rect 4566 4868 4570 4924
rect 4506 4864 4570 4868
rect 4586 4924 4650 4928
rect 4586 4868 4590 4924
rect 4590 4868 4646 4924
rect 4646 4868 4650 4924
rect 4586 4864 4650 4868
rect 4666 4924 4730 4928
rect 4666 4868 4670 4924
rect 4670 4868 4726 4924
rect 4726 4868 4730 4924
rect 4666 4864 4730 4868
rect 11374 4924 11438 4928
rect 11374 4868 11378 4924
rect 11378 4868 11434 4924
rect 11434 4868 11438 4924
rect 11374 4864 11438 4868
rect 11454 4924 11518 4928
rect 11454 4868 11458 4924
rect 11458 4868 11514 4924
rect 11514 4868 11518 4924
rect 11454 4864 11518 4868
rect 11534 4924 11598 4928
rect 11534 4868 11538 4924
rect 11538 4868 11594 4924
rect 11594 4868 11598 4924
rect 11534 4864 11598 4868
rect 11614 4924 11678 4928
rect 11614 4868 11618 4924
rect 11618 4868 11674 4924
rect 11674 4868 11678 4924
rect 11614 4864 11678 4868
rect 18322 4924 18386 4928
rect 18322 4868 18326 4924
rect 18326 4868 18382 4924
rect 18382 4868 18386 4924
rect 18322 4864 18386 4868
rect 18402 4924 18466 4928
rect 18402 4868 18406 4924
rect 18406 4868 18462 4924
rect 18462 4868 18466 4924
rect 18402 4864 18466 4868
rect 18482 4924 18546 4928
rect 18482 4868 18486 4924
rect 18486 4868 18542 4924
rect 18542 4868 18546 4924
rect 18482 4864 18546 4868
rect 18562 4924 18626 4928
rect 18562 4868 18566 4924
rect 18566 4868 18622 4924
rect 18622 4868 18626 4924
rect 18562 4864 18626 4868
rect 25270 4924 25334 4928
rect 25270 4868 25274 4924
rect 25274 4868 25330 4924
rect 25330 4868 25334 4924
rect 25270 4864 25334 4868
rect 25350 4924 25414 4928
rect 25350 4868 25354 4924
rect 25354 4868 25410 4924
rect 25410 4868 25414 4924
rect 25350 4864 25414 4868
rect 25430 4924 25494 4928
rect 25430 4868 25434 4924
rect 25434 4868 25490 4924
rect 25490 4868 25494 4924
rect 25430 4864 25494 4868
rect 25510 4924 25574 4928
rect 25510 4868 25514 4924
rect 25514 4868 25570 4924
rect 25570 4868 25574 4924
rect 25510 4864 25574 4868
rect 7900 4380 7964 4384
rect 7900 4324 7904 4380
rect 7904 4324 7960 4380
rect 7960 4324 7964 4380
rect 7900 4320 7964 4324
rect 7980 4380 8044 4384
rect 7980 4324 7984 4380
rect 7984 4324 8040 4380
rect 8040 4324 8044 4380
rect 7980 4320 8044 4324
rect 8060 4380 8124 4384
rect 8060 4324 8064 4380
rect 8064 4324 8120 4380
rect 8120 4324 8124 4380
rect 8060 4320 8124 4324
rect 8140 4380 8204 4384
rect 8140 4324 8144 4380
rect 8144 4324 8200 4380
rect 8200 4324 8204 4380
rect 8140 4320 8204 4324
rect 14848 4380 14912 4384
rect 14848 4324 14852 4380
rect 14852 4324 14908 4380
rect 14908 4324 14912 4380
rect 14848 4320 14912 4324
rect 14928 4380 14992 4384
rect 14928 4324 14932 4380
rect 14932 4324 14988 4380
rect 14988 4324 14992 4380
rect 14928 4320 14992 4324
rect 15008 4380 15072 4384
rect 15008 4324 15012 4380
rect 15012 4324 15068 4380
rect 15068 4324 15072 4380
rect 15008 4320 15072 4324
rect 15088 4380 15152 4384
rect 15088 4324 15092 4380
rect 15092 4324 15148 4380
rect 15148 4324 15152 4380
rect 15088 4320 15152 4324
rect 21796 4380 21860 4384
rect 21796 4324 21800 4380
rect 21800 4324 21856 4380
rect 21856 4324 21860 4380
rect 21796 4320 21860 4324
rect 21876 4380 21940 4384
rect 21876 4324 21880 4380
rect 21880 4324 21936 4380
rect 21936 4324 21940 4380
rect 21876 4320 21940 4324
rect 21956 4380 22020 4384
rect 21956 4324 21960 4380
rect 21960 4324 22016 4380
rect 22016 4324 22020 4380
rect 21956 4320 22020 4324
rect 22036 4380 22100 4384
rect 22036 4324 22040 4380
rect 22040 4324 22096 4380
rect 22096 4324 22100 4380
rect 22036 4320 22100 4324
rect 4426 3836 4490 3840
rect 4426 3780 4430 3836
rect 4430 3780 4486 3836
rect 4486 3780 4490 3836
rect 4426 3776 4490 3780
rect 4506 3836 4570 3840
rect 4506 3780 4510 3836
rect 4510 3780 4566 3836
rect 4566 3780 4570 3836
rect 4506 3776 4570 3780
rect 4586 3836 4650 3840
rect 4586 3780 4590 3836
rect 4590 3780 4646 3836
rect 4646 3780 4650 3836
rect 4586 3776 4650 3780
rect 4666 3836 4730 3840
rect 4666 3780 4670 3836
rect 4670 3780 4726 3836
rect 4726 3780 4730 3836
rect 4666 3776 4730 3780
rect 11374 3836 11438 3840
rect 11374 3780 11378 3836
rect 11378 3780 11434 3836
rect 11434 3780 11438 3836
rect 11374 3776 11438 3780
rect 11454 3836 11518 3840
rect 11454 3780 11458 3836
rect 11458 3780 11514 3836
rect 11514 3780 11518 3836
rect 11454 3776 11518 3780
rect 11534 3836 11598 3840
rect 11534 3780 11538 3836
rect 11538 3780 11594 3836
rect 11594 3780 11598 3836
rect 11534 3776 11598 3780
rect 11614 3836 11678 3840
rect 11614 3780 11618 3836
rect 11618 3780 11674 3836
rect 11674 3780 11678 3836
rect 11614 3776 11678 3780
rect 18322 3836 18386 3840
rect 18322 3780 18326 3836
rect 18326 3780 18382 3836
rect 18382 3780 18386 3836
rect 18322 3776 18386 3780
rect 18402 3836 18466 3840
rect 18402 3780 18406 3836
rect 18406 3780 18462 3836
rect 18462 3780 18466 3836
rect 18402 3776 18466 3780
rect 18482 3836 18546 3840
rect 18482 3780 18486 3836
rect 18486 3780 18542 3836
rect 18542 3780 18546 3836
rect 18482 3776 18546 3780
rect 18562 3836 18626 3840
rect 18562 3780 18566 3836
rect 18566 3780 18622 3836
rect 18622 3780 18626 3836
rect 18562 3776 18626 3780
rect 25270 3836 25334 3840
rect 25270 3780 25274 3836
rect 25274 3780 25330 3836
rect 25330 3780 25334 3836
rect 25270 3776 25334 3780
rect 25350 3836 25414 3840
rect 25350 3780 25354 3836
rect 25354 3780 25410 3836
rect 25410 3780 25414 3836
rect 25350 3776 25414 3780
rect 25430 3836 25494 3840
rect 25430 3780 25434 3836
rect 25434 3780 25490 3836
rect 25490 3780 25494 3836
rect 25430 3776 25494 3780
rect 25510 3836 25574 3840
rect 25510 3780 25514 3836
rect 25514 3780 25570 3836
rect 25570 3780 25574 3836
rect 25510 3776 25574 3780
rect 7900 3292 7964 3296
rect 7900 3236 7904 3292
rect 7904 3236 7960 3292
rect 7960 3236 7964 3292
rect 7900 3232 7964 3236
rect 7980 3292 8044 3296
rect 7980 3236 7984 3292
rect 7984 3236 8040 3292
rect 8040 3236 8044 3292
rect 7980 3232 8044 3236
rect 8060 3292 8124 3296
rect 8060 3236 8064 3292
rect 8064 3236 8120 3292
rect 8120 3236 8124 3292
rect 8060 3232 8124 3236
rect 8140 3292 8204 3296
rect 8140 3236 8144 3292
rect 8144 3236 8200 3292
rect 8200 3236 8204 3292
rect 8140 3232 8204 3236
rect 14848 3292 14912 3296
rect 14848 3236 14852 3292
rect 14852 3236 14908 3292
rect 14908 3236 14912 3292
rect 14848 3232 14912 3236
rect 14928 3292 14992 3296
rect 14928 3236 14932 3292
rect 14932 3236 14988 3292
rect 14988 3236 14992 3292
rect 14928 3232 14992 3236
rect 15008 3292 15072 3296
rect 15008 3236 15012 3292
rect 15012 3236 15068 3292
rect 15068 3236 15072 3292
rect 15008 3232 15072 3236
rect 15088 3292 15152 3296
rect 15088 3236 15092 3292
rect 15092 3236 15148 3292
rect 15148 3236 15152 3292
rect 15088 3232 15152 3236
rect 21796 3292 21860 3296
rect 21796 3236 21800 3292
rect 21800 3236 21856 3292
rect 21856 3236 21860 3292
rect 21796 3232 21860 3236
rect 21876 3292 21940 3296
rect 21876 3236 21880 3292
rect 21880 3236 21936 3292
rect 21936 3236 21940 3292
rect 21876 3232 21940 3236
rect 21956 3292 22020 3296
rect 21956 3236 21960 3292
rect 21960 3236 22016 3292
rect 22016 3236 22020 3292
rect 21956 3232 22020 3236
rect 22036 3292 22100 3296
rect 22036 3236 22040 3292
rect 22040 3236 22096 3292
rect 22096 3236 22100 3292
rect 22036 3232 22100 3236
rect 4426 2748 4490 2752
rect 4426 2692 4430 2748
rect 4430 2692 4486 2748
rect 4486 2692 4490 2748
rect 4426 2688 4490 2692
rect 4506 2748 4570 2752
rect 4506 2692 4510 2748
rect 4510 2692 4566 2748
rect 4566 2692 4570 2748
rect 4506 2688 4570 2692
rect 4586 2748 4650 2752
rect 4586 2692 4590 2748
rect 4590 2692 4646 2748
rect 4646 2692 4650 2748
rect 4586 2688 4650 2692
rect 4666 2748 4730 2752
rect 4666 2692 4670 2748
rect 4670 2692 4726 2748
rect 4726 2692 4730 2748
rect 4666 2688 4730 2692
rect 11374 2748 11438 2752
rect 11374 2692 11378 2748
rect 11378 2692 11434 2748
rect 11434 2692 11438 2748
rect 11374 2688 11438 2692
rect 11454 2748 11518 2752
rect 11454 2692 11458 2748
rect 11458 2692 11514 2748
rect 11514 2692 11518 2748
rect 11454 2688 11518 2692
rect 11534 2748 11598 2752
rect 11534 2692 11538 2748
rect 11538 2692 11594 2748
rect 11594 2692 11598 2748
rect 11534 2688 11598 2692
rect 11614 2748 11678 2752
rect 11614 2692 11618 2748
rect 11618 2692 11674 2748
rect 11674 2692 11678 2748
rect 11614 2688 11678 2692
rect 18322 2748 18386 2752
rect 18322 2692 18326 2748
rect 18326 2692 18382 2748
rect 18382 2692 18386 2748
rect 18322 2688 18386 2692
rect 18402 2748 18466 2752
rect 18402 2692 18406 2748
rect 18406 2692 18462 2748
rect 18462 2692 18466 2748
rect 18402 2688 18466 2692
rect 18482 2748 18546 2752
rect 18482 2692 18486 2748
rect 18486 2692 18542 2748
rect 18542 2692 18546 2748
rect 18482 2688 18546 2692
rect 18562 2748 18626 2752
rect 18562 2692 18566 2748
rect 18566 2692 18622 2748
rect 18622 2692 18626 2748
rect 18562 2688 18626 2692
rect 25270 2748 25334 2752
rect 25270 2692 25274 2748
rect 25274 2692 25330 2748
rect 25330 2692 25334 2748
rect 25270 2688 25334 2692
rect 25350 2748 25414 2752
rect 25350 2692 25354 2748
rect 25354 2692 25410 2748
rect 25410 2692 25414 2748
rect 25350 2688 25414 2692
rect 25430 2748 25494 2752
rect 25430 2692 25434 2748
rect 25434 2692 25490 2748
rect 25490 2692 25494 2748
rect 25430 2688 25494 2692
rect 25510 2748 25574 2752
rect 25510 2692 25514 2748
rect 25514 2692 25570 2748
rect 25570 2692 25574 2748
rect 25510 2688 25574 2692
rect 7900 2204 7964 2208
rect 7900 2148 7904 2204
rect 7904 2148 7960 2204
rect 7960 2148 7964 2204
rect 7900 2144 7964 2148
rect 7980 2204 8044 2208
rect 7980 2148 7984 2204
rect 7984 2148 8040 2204
rect 8040 2148 8044 2204
rect 7980 2144 8044 2148
rect 8060 2204 8124 2208
rect 8060 2148 8064 2204
rect 8064 2148 8120 2204
rect 8120 2148 8124 2204
rect 8060 2144 8124 2148
rect 8140 2204 8204 2208
rect 8140 2148 8144 2204
rect 8144 2148 8200 2204
rect 8200 2148 8204 2204
rect 8140 2144 8204 2148
rect 14848 2204 14912 2208
rect 14848 2148 14852 2204
rect 14852 2148 14908 2204
rect 14908 2148 14912 2204
rect 14848 2144 14912 2148
rect 14928 2204 14992 2208
rect 14928 2148 14932 2204
rect 14932 2148 14988 2204
rect 14988 2148 14992 2204
rect 14928 2144 14992 2148
rect 15008 2204 15072 2208
rect 15008 2148 15012 2204
rect 15012 2148 15068 2204
rect 15068 2148 15072 2204
rect 15008 2144 15072 2148
rect 15088 2204 15152 2208
rect 15088 2148 15092 2204
rect 15092 2148 15148 2204
rect 15148 2148 15152 2204
rect 15088 2144 15152 2148
rect 21796 2204 21860 2208
rect 21796 2148 21800 2204
rect 21800 2148 21856 2204
rect 21856 2148 21860 2204
rect 21796 2144 21860 2148
rect 21876 2204 21940 2208
rect 21876 2148 21880 2204
rect 21880 2148 21936 2204
rect 21936 2148 21940 2204
rect 21876 2144 21940 2148
rect 21956 2204 22020 2208
rect 21956 2148 21960 2204
rect 21960 2148 22016 2204
rect 22016 2148 22020 2204
rect 21956 2144 22020 2148
rect 22036 2204 22100 2208
rect 22036 2148 22040 2204
rect 22040 2148 22096 2204
rect 22096 2148 22100 2204
rect 22036 2144 22100 2148
<< metal4 >>
rect 4418 27776 4738 27792
rect 4418 27712 4426 27776
rect 4490 27712 4506 27776
rect 4570 27712 4586 27776
rect 4650 27712 4666 27776
rect 4730 27712 4738 27776
rect 4418 26688 4738 27712
rect 4418 26624 4426 26688
rect 4490 26624 4506 26688
rect 4570 26624 4586 26688
rect 4650 26624 4666 26688
rect 4730 26624 4738 26688
rect 4418 25600 4738 26624
rect 4418 25536 4426 25600
rect 4490 25536 4506 25600
rect 4570 25536 4586 25600
rect 4650 25536 4666 25600
rect 4730 25536 4738 25600
rect 4418 24512 4738 25536
rect 4418 24448 4426 24512
rect 4490 24448 4506 24512
rect 4570 24448 4586 24512
rect 4650 24448 4666 24512
rect 4730 24448 4738 24512
rect 4418 23424 4738 24448
rect 4418 23360 4426 23424
rect 4490 23360 4506 23424
rect 4570 23360 4586 23424
rect 4650 23360 4666 23424
rect 4730 23360 4738 23424
rect 4418 22336 4738 23360
rect 4418 22272 4426 22336
rect 4490 22272 4506 22336
rect 4570 22272 4586 22336
rect 4650 22272 4666 22336
rect 4730 22272 4738 22336
rect 4418 21248 4738 22272
rect 4418 21184 4426 21248
rect 4490 21184 4506 21248
rect 4570 21184 4586 21248
rect 4650 21184 4666 21248
rect 4730 21184 4738 21248
rect 4418 20160 4738 21184
rect 4418 20096 4426 20160
rect 4490 20096 4506 20160
rect 4570 20096 4586 20160
rect 4650 20096 4666 20160
rect 4730 20096 4738 20160
rect 4418 19072 4738 20096
rect 4418 19008 4426 19072
rect 4490 19008 4506 19072
rect 4570 19008 4586 19072
rect 4650 19008 4666 19072
rect 4730 19008 4738 19072
rect 4418 17984 4738 19008
rect 4418 17920 4426 17984
rect 4490 17920 4506 17984
rect 4570 17920 4586 17984
rect 4650 17920 4666 17984
rect 4730 17920 4738 17984
rect 4418 16896 4738 17920
rect 4418 16832 4426 16896
rect 4490 16832 4506 16896
rect 4570 16832 4586 16896
rect 4650 16832 4666 16896
rect 4730 16832 4738 16896
rect 4418 15808 4738 16832
rect 4418 15744 4426 15808
rect 4490 15744 4506 15808
rect 4570 15744 4586 15808
rect 4650 15744 4666 15808
rect 4730 15744 4738 15808
rect 4418 14720 4738 15744
rect 4418 14656 4426 14720
rect 4490 14656 4506 14720
rect 4570 14656 4586 14720
rect 4650 14656 4666 14720
rect 4730 14656 4738 14720
rect 4418 13632 4738 14656
rect 4418 13568 4426 13632
rect 4490 13568 4506 13632
rect 4570 13568 4586 13632
rect 4650 13568 4666 13632
rect 4730 13568 4738 13632
rect 4418 12544 4738 13568
rect 4418 12480 4426 12544
rect 4490 12480 4506 12544
rect 4570 12480 4586 12544
rect 4650 12480 4666 12544
rect 4730 12480 4738 12544
rect 4418 11456 4738 12480
rect 4418 11392 4426 11456
rect 4490 11392 4506 11456
rect 4570 11392 4586 11456
rect 4650 11392 4666 11456
rect 4730 11392 4738 11456
rect 4418 10368 4738 11392
rect 4418 10304 4426 10368
rect 4490 10304 4506 10368
rect 4570 10304 4586 10368
rect 4650 10304 4666 10368
rect 4730 10304 4738 10368
rect 4418 9280 4738 10304
rect 4418 9216 4426 9280
rect 4490 9216 4506 9280
rect 4570 9216 4586 9280
rect 4650 9216 4666 9280
rect 4730 9216 4738 9280
rect 4418 8192 4738 9216
rect 4418 8128 4426 8192
rect 4490 8128 4506 8192
rect 4570 8128 4586 8192
rect 4650 8128 4666 8192
rect 4730 8128 4738 8192
rect 4418 7104 4738 8128
rect 4418 7040 4426 7104
rect 4490 7040 4506 7104
rect 4570 7040 4586 7104
rect 4650 7040 4666 7104
rect 4730 7040 4738 7104
rect 4418 6016 4738 7040
rect 4418 5952 4426 6016
rect 4490 5952 4506 6016
rect 4570 5952 4586 6016
rect 4650 5952 4666 6016
rect 4730 5952 4738 6016
rect 4418 4928 4738 5952
rect 4418 4864 4426 4928
rect 4490 4864 4506 4928
rect 4570 4864 4586 4928
rect 4650 4864 4666 4928
rect 4730 4864 4738 4928
rect 4418 3840 4738 4864
rect 4418 3776 4426 3840
rect 4490 3776 4506 3840
rect 4570 3776 4586 3840
rect 4650 3776 4666 3840
rect 4730 3776 4738 3840
rect 4418 2752 4738 3776
rect 4418 2688 4426 2752
rect 4490 2688 4506 2752
rect 4570 2688 4586 2752
rect 4650 2688 4666 2752
rect 4730 2688 4738 2752
rect 4418 2128 4738 2688
rect 7892 27232 8212 27792
rect 7892 27168 7900 27232
rect 7964 27168 7980 27232
rect 8044 27168 8060 27232
rect 8124 27168 8140 27232
rect 8204 27168 8212 27232
rect 7892 26144 8212 27168
rect 7892 26080 7900 26144
rect 7964 26080 7980 26144
rect 8044 26080 8060 26144
rect 8124 26080 8140 26144
rect 8204 26080 8212 26144
rect 7892 25056 8212 26080
rect 7892 24992 7900 25056
rect 7964 24992 7980 25056
rect 8044 24992 8060 25056
rect 8124 24992 8140 25056
rect 8204 24992 8212 25056
rect 7892 23968 8212 24992
rect 7892 23904 7900 23968
rect 7964 23904 7980 23968
rect 8044 23904 8060 23968
rect 8124 23904 8140 23968
rect 8204 23904 8212 23968
rect 7892 22880 8212 23904
rect 7892 22816 7900 22880
rect 7964 22816 7980 22880
rect 8044 22816 8060 22880
rect 8124 22816 8140 22880
rect 8204 22816 8212 22880
rect 7892 21792 8212 22816
rect 7892 21728 7900 21792
rect 7964 21728 7980 21792
rect 8044 21728 8060 21792
rect 8124 21728 8140 21792
rect 8204 21728 8212 21792
rect 7892 20704 8212 21728
rect 7892 20640 7900 20704
rect 7964 20640 7980 20704
rect 8044 20640 8060 20704
rect 8124 20640 8140 20704
rect 8204 20640 8212 20704
rect 7892 19616 8212 20640
rect 7892 19552 7900 19616
rect 7964 19552 7980 19616
rect 8044 19552 8060 19616
rect 8124 19552 8140 19616
rect 8204 19552 8212 19616
rect 7892 18528 8212 19552
rect 7892 18464 7900 18528
rect 7964 18464 7980 18528
rect 8044 18464 8060 18528
rect 8124 18464 8140 18528
rect 8204 18464 8212 18528
rect 7892 17440 8212 18464
rect 7892 17376 7900 17440
rect 7964 17376 7980 17440
rect 8044 17376 8060 17440
rect 8124 17376 8140 17440
rect 8204 17376 8212 17440
rect 7892 16352 8212 17376
rect 7892 16288 7900 16352
rect 7964 16288 7980 16352
rect 8044 16288 8060 16352
rect 8124 16288 8140 16352
rect 8204 16288 8212 16352
rect 7892 15264 8212 16288
rect 7892 15200 7900 15264
rect 7964 15200 7980 15264
rect 8044 15200 8060 15264
rect 8124 15200 8140 15264
rect 8204 15200 8212 15264
rect 7892 14176 8212 15200
rect 7892 14112 7900 14176
rect 7964 14112 7980 14176
rect 8044 14112 8060 14176
rect 8124 14112 8140 14176
rect 8204 14112 8212 14176
rect 7892 13088 8212 14112
rect 7892 13024 7900 13088
rect 7964 13024 7980 13088
rect 8044 13024 8060 13088
rect 8124 13024 8140 13088
rect 8204 13024 8212 13088
rect 7892 12000 8212 13024
rect 7892 11936 7900 12000
rect 7964 11936 7980 12000
rect 8044 11936 8060 12000
rect 8124 11936 8140 12000
rect 8204 11936 8212 12000
rect 7892 10912 8212 11936
rect 7892 10848 7900 10912
rect 7964 10848 7980 10912
rect 8044 10848 8060 10912
rect 8124 10848 8140 10912
rect 8204 10848 8212 10912
rect 7892 9824 8212 10848
rect 7892 9760 7900 9824
rect 7964 9760 7980 9824
rect 8044 9760 8060 9824
rect 8124 9760 8140 9824
rect 8204 9760 8212 9824
rect 7892 8736 8212 9760
rect 7892 8672 7900 8736
rect 7964 8672 7980 8736
rect 8044 8672 8060 8736
rect 8124 8672 8140 8736
rect 8204 8672 8212 8736
rect 7892 7648 8212 8672
rect 7892 7584 7900 7648
rect 7964 7584 7980 7648
rect 8044 7584 8060 7648
rect 8124 7584 8140 7648
rect 8204 7584 8212 7648
rect 7892 6560 8212 7584
rect 7892 6496 7900 6560
rect 7964 6496 7980 6560
rect 8044 6496 8060 6560
rect 8124 6496 8140 6560
rect 8204 6496 8212 6560
rect 7892 5472 8212 6496
rect 7892 5408 7900 5472
rect 7964 5408 7980 5472
rect 8044 5408 8060 5472
rect 8124 5408 8140 5472
rect 8204 5408 8212 5472
rect 7892 4384 8212 5408
rect 7892 4320 7900 4384
rect 7964 4320 7980 4384
rect 8044 4320 8060 4384
rect 8124 4320 8140 4384
rect 8204 4320 8212 4384
rect 7892 3296 8212 4320
rect 7892 3232 7900 3296
rect 7964 3232 7980 3296
rect 8044 3232 8060 3296
rect 8124 3232 8140 3296
rect 8204 3232 8212 3296
rect 7892 2208 8212 3232
rect 7892 2144 7900 2208
rect 7964 2144 7980 2208
rect 8044 2144 8060 2208
rect 8124 2144 8140 2208
rect 8204 2144 8212 2208
rect 7892 2128 8212 2144
rect 11366 27776 11686 27792
rect 11366 27712 11374 27776
rect 11438 27712 11454 27776
rect 11518 27712 11534 27776
rect 11598 27712 11614 27776
rect 11678 27712 11686 27776
rect 11366 26688 11686 27712
rect 11366 26624 11374 26688
rect 11438 26624 11454 26688
rect 11518 26624 11534 26688
rect 11598 26624 11614 26688
rect 11678 26624 11686 26688
rect 11366 25600 11686 26624
rect 11366 25536 11374 25600
rect 11438 25536 11454 25600
rect 11518 25536 11534 25600
rect 11598 25536 11614 25600
rect 11678 25536 11686 25600
rect 11366 24512 11686 25536
rect 11366 24448 11374 24512
rect 11438 24448 11454 24512
rect 11518 24448 11534 24512
rect 11598 24448 11614 24512
rect 11678 24448 11686 24512
rect 11366 23424 11686 24448
rect 11366 23360 11374 23424
rect 11438 23360 11454 23424
rect 11518 23360 11534 23424
rect 11598 23360 11614 23424
rect 11678 23360 11686 23424
rect 11366 22336 11686 23360
rect 11366 22272 11374 22336
rect 11438 22272 11454 22336
rect 11518 22272 11534 22336
rect 11598 22272 11614 22336
rect 11678 22272 11686 22336
rect 11366 21248 11686 22272
rect 11366 21184 11374 21248
rect 11438 21184 11454 21248
rect 11518 21184 11534 21248
rect 11598 21184 11614 21248
rect 11678 21184 11686 21248
rect 11366 20160 11686 21184
rect 11366 20096 11374 20160
rect 11438 20096 11454 20160
rect 11518 20096 11534 20160
rect 11598 20096 11614 20160
rect 11678 20096 11686 20160
rect 11366 19072 11686 20096
rect 11366 19008 11374 19072
rect 11438 19008 11454 19072
rect 11518 19008 11534 19072
rect 11598 19008 11614 19072
rect 11678 19008 11686 19072
rect 11366 17984 11686 19008
rect 11366 17920 11374 17984
rect 11438 17920 11454 17984
rect 11518 17920 11534 17984
rect 11598 17920 11614 17984
rect 11678 17920 11686 17984
rect 11366 16896 11686 17920
rect 11366 16832 11374 16896
rect 11438 16832 11454 16896
rect 11518 16832 11534 16896
rect 11598 16832 11614 16896
rect 11678 16832 11686 16896
rect 11366 15808 11686 16832
rect 11366 15744 11374 15808
rect 11438 15744 11454 15808
rect 11518 15744 11534 15808
rect 11598 15744 11614 15808
rect 11678 15744 11686 15808
rect 11366 14720 11686 15744
rect 11366 14656 11374 14720
rect 11438 14656 11454 14720
rect 11518 14656 11534 14720
rect 11598 14656 11614 14720
rect 11678 14656 11686 14720
rect 11366 13632 11686 14656
rect 11366 13568 11374 13632
rect 11438 13568 11454 13632
rect 11518 13568 11534 13632
rect 11598 13568 11614 13632
rect 11678 13568 11686 13632
rect 11366 12544 11686 13568
rect 11366 12480 11374 12544
rect 11438 12480 11454 12544
rect 11518 12480 11534 12544
rect 11598 12480 11614 12544
rect 11678 12480 11686 12544
rect 11366 11456 11686 12480
rect 11366 11392 11374 11456
rect 11438 11392 11454 11456
rect 11518 11392 11534 11456
rect 11598 11392 11614 11456
rect 11678 11392 11686 11456
rect 11366 10368 11686 11392
rect 11366 10304 11374 10368
rect 11438 10304 11454 10368
rect 11518 10304 11534 10368
rect 11598 10304 11614 10368
rect 11678 10304 11686 10368
rect 11366 9280 11686 10304
rect 11366 9216 11374 9280
rect 11438 9216 11454 9280
rect 11518 9216 11534 9280
rect 11598 9216 11614 9280
rect 11678 9216 11686 9280
rect 11366 8192 11686 9216
rect 11366 8128 11374 8192
rect 11438 8128 11454 8192
rect 11518 8128 11534 8192
rect 11598 8128 11614 8192
rect 11678 8128 11686 8192
rect 11366 7104 11686 8128
rect 11366 7040 11374 7104
rect 11438 7040 11454 7104
rect 11518 7040 11534 7104
rect 11598 7040 11614 7104
rect 11678 7040 11686 7104
rect 11366 6016 11686 7040
rect 11366 5952 11374 6016
rect 11438 5952 11454 6016
rect 11518 5952 11534 6016
rect 11598 5952 11614 6016
rect 11678 5952 11686 6016
rect 11366 4928 11686 5952
rect 11366 4864 11374 4928
rect 11438 4864 11454 4928
rect 11518 4864 11534 4928
rect 11598 4864 11614 4928
rect 11678 4864 11686 4928
rect 11366 3840 11686 4864
rect 11366 3776 11374 3840
rect 11438 3776 11454 3840
rect 11518 3776 11534 3840
rect 11598 3776 11614 3840
rect 11678 3776 11686 3840
rect 11366 2752 11686 3776
rect 11366 2688 11374 2752
rect 11438 2688 11454 2752
rect 11518 2688 11534 2752
rect 11598 2688 11614 2752
rect 11678 2688 11686 2752
rect 11366 2128 11686 2688
rect 14840 27232 15160 27792
rect 14840 27168 14848 27232
rect 14912 27168 14928 27232
rect 14992 27168 15008 27232
rect 15072 27168 15088 27232
rect 15152 27168 15160 27232
rect 14840 26144 15160 27168
rect 14840 26080 14848 26144
rect 14912 26080 14928 26144
rect 14992 26080 15008 26144
rect 15072 26080 15088 26144
rect 15152 26080 15160 26144
rect 14840 25056 15160 26080
rect 14840 24992 14848 25056
rect 14912 24992 14928 25056
rect 14992 24992 15008 25056
rect 15072 24992 15088 25056
rect 15152 24992 15160 25056
rect 14840 23968 15160 24992
rect 14840 23904 14848 23968
rect 14912 23904 14928 23968
rect 14992 23904 15008 23968
rect 15072 23904 15088 23968
rect 15152 23904 15160 23968
rect 14840 22880 15160 23904
rect 14840 22816 14848 22880
rect 14912 22816 14928 22880
rect 14992 22816 15008 22880
rect 15072 22816 15088 22880
rect 15152 22816 15160 22880
rect 14840 21792 15160 22816
rect 14840 21728 14848 21792
rect 14912 21728 14928 21792
rect 14992 21728 15008 21792
rect 15072 21728 15088 21792
rect 15152 21728 15160 21792
rect 14840 20704 15160 21728
rect 14840 20640 14848 20704
rect 14912 20640 14928 20704
rect 14992 20640 15008 20704
rect 15072 20640 15088 20704
rect 15152 20640 15160 20704
rect 14840 19616 15160 20640
rect 14840 19552 14848 19616
rect 14912 19552 14928 19616
rect 14992 19552 15008 19616
rect 15072 19552 15088 19616
rect 15152 19552 15160 19616
rect 14840 18528 15160 19552
rect 14840 18464 14848 18528
rect 14912 18464 14928 18528
rect 14992 18464 15008 18528
rect 15072 18464 15088 18528
rect 15152 18464 15160 18528
rect 14840 17440 15160 18464
rect 14840 17376 14848 17440
rect 14912 17376 14928 17440
rect 14992 17376 15008 17440
rect 15072 17376 15088 17440
rect 15152 17376 15160 17440
rect 14840 16352 15160 17376
rect 14840 16288 14848 16352
rect 14912 16288 14928 16352
rect 14992 16288 15008 16352
rect 15072 16288 15088 16352
rect 15152 16288 15160 16352
rect 14840 15264 15160 16288
rect 14840 15200 14848 15264
rect 14912 15200 14928 15264
rect 14992 15200 15008 15264
rect 15072 15200 15088 15264
rect 15152 15200 15160 15264
rect 14840 14176 15160 15200
rect 14840 14112 14848 14176
rect 14912 14112 14928 14176
rect 14992 14112 15008 14176
rect 15072 14112 15088 14176
rect 15152 14112 15160 14176
rect 14840 13088 15160 14112
rect 14840 13024 14848 13088
rect 14912 13024 14928 13088
rect 14992 13024 15008 13088
rect 15072 13024 15088 13088
rect 15152 13024 15160 13088
rect 14840 12000 15160 13024
rect 14840 11936 14848 12000
rect 14912 11936 14928 12000
rect 14992 11936 15008 12000
rect 15072 11936 15088 12000
rect 15152 11936 15160 12000
rect 14840 10912 15160 11936
rect 14840 10848 14848 10912
rect 14912 10848 14928 10912
rect 14992 10848 15008 10912
rect 15072 10848 15088 10912
rect 15152 10848 15160 10912
rect 14840 9824 15160 10848
rect 14840 9760 14848 9824
rect 14912 9760 14928 9824
rect 14992 9760 15008 9824
rect 15072 9760 15088 9824
rect 15152 9760 15160 9824
rect 14840 8736 15160 9760
rect 14840 8672 14848 8736
rect 14912 8672 14928 8736
rect 14992 8672 15008 8736
rect 15072 8672 15088 8736
rect 15152 8672 15160 8736
rect 14840 7648 15160 8672
rect 14840 7584 14848 7648
rect 14912 7584 14928 7648
rect 14992 7584 15008 7648
rect 15072 7584 15088 7648
rect 15152 7584 15160 7648
rect 14840 6560 15160 7584
rect 14840 6496 14848 6560
rect 14912 6496 14928 6560
rect 14992 6496 15008 6560
rect 15072 6496 15088 6560
rect 15152 6496 15160 6560
rect 14840 5472 15160 6496
rect 14840 5408 14848 5472
rect 14912 5408 14928 5472
rect 14992 5408 15008 5472
rect 15072 5408 15088 5472
rect 15152 5408 15160 5472
rect 14840 4384 15160 5408
rect 14840 4320 14848 4384
rect 14912 4320 14928 4384
rect 14992 4320 15008 4384
rect 15072 4320 15088 4384
rect 15152 4320 15160 4384
rect 14840 3296 15160 4320
rect 14840 3232 14848 3296
rect 14912 3232 14928 3296
rect 14992 3232 15008 3296
rect 15072 3232 15088 3296
rect 15152 3232 15160 3296
rect 14840 2208 15160 3232
rect 14840 2144 14848 2208
rect 14912 2144 14928 2208
rect 14992 2144 15008 2208
rect 15072 2144 15088 2208
rect 15152 2144 15160 2208
rect 14840 2128 15160 2144
rect 18314 27776 18634 27792
rect 18314 27712 18322 27776
rect 18386 27712 18402 27776
rect 18466 27712 18482 27776
rect 18546 27712 18562 27776
rect 18626 27712 18634 27776
rect 18314 26688 18634 27712
rect 18314 26624 18322 26688
rect 18386 26624 18402 26688
rect 18466 26624 18482 26688
rect 18546 26624 18562 26688
rect 18626 26624 18634 26688
rect 18314 25600 18634 26624
rect 18314 25536 18322 25600
rect 18386 25536 18402 25600
rect 18466 25536 18482 25600
rect 18546 25536 18562 25600
rect 18626 25536 18634 25600
rect 18314 24512 18634 25536
rect 18314 24448 18322 24512
rect 18386 24448 18402 24512
rect 18466 24448 18482 24512
rect 18546 24448 18562 24512
rect 18626 24448 18634 24512
rect 18314 23424 18634 24448
rect 18314 23360 18322 23424
rect 18386 23360 18402 23424
rect 18466 23360 18482 23424
rect 18546 23360 18562 23424
rect 18626 23360 18634 23424
rect 18314 22336 18634 23360
rect 18314 22272 18322 22336
rect 18386 22272 18402 22336
rect 18466 22272 18482 22336
rect 18546 22272 18562 22336
rect 18626 22272 18634 22336
rect 18314 21248 18634 22272
rect 18314 21184 18322 21248
rect 18386 21184 18402 21248
rect 18466 21184 18482 21248
rect 18546 21184 18562 21248
rect 18626 21184 18634 21248
rect 18314 20160 18634 21184
rect 18314 20096 18322 20160
rect 18386 20096 18402 20160
rect 18466 20096 18482 20160
rect 18546 20096 18562 20160
rect 18626 20096 18634 20160
rect 18314 19072 18634 20096
rect 18314 19008 18322 19072
rect 18386 19008 18402 19072
rect 18466 19008 18482 19072
rect 18546 19008 18562 19072
rect 18626 19008 18634 19072
rect 18314 17984 18634 19008
rect 18314 17920 18322 17984
rect 18386 17920 18402 17984
rect 18466 17920 18482 17984
rect 18546 17920 18562 17984
rect 18626 17920 18634 17984
rect 18314 16896 18634 17920
rect 18314 16832 18322 16896
rect 18386 16832 18402 16896
rect 18466 16832 18482 16896
rect 18546 16832 18562 16896
rect 18626 16832 18634 16896
rect 18314 15808 18634 16832
rect 18314 15744 18322 15808
rect 18386 15744 18402 15808
rect 18466 15744 18482 15808
rect 18546 15744 18562 15808
rect 18626 15744 18634 15808
rect 18314 14720 18634 15744
rect 18314 14656 18322 14720
rect 18386 14656 18402 14720
rect 18466 14656 18482 14720
rect 18546 14656 18562 14720
rect 18626 14656 18634 14720
rect 18314 13632 18634 14656
rect 18314 13568 18322 13632
rect 18386 13568 18402 13632
rect 18466 13568 18482 13632
rect 18546 13568 18562 13632
rect 18626 13568 18634 13632
rect 18314 12544 18634 13568
rect 18314 12480 18322 12544
rect 18386 12480 18402 12544
rect 18466 12480 18482 12544
rect 18546 12480 18562 12544
rect 18626 12480 18634 12544
rect 18314 11456 18634 12480
rect 18314 11392 18322 11456
rect 18386 11392 18402 11456
rect 18466 11392 18482 11456
rect 18546 11392 18562 11456
rect 18626 11392 18634 11456
rect 18314 10368 18634 11392
rect 18314 10304 18322 10368
rect 18386 10304 18402 10368
rect 18466 10304 18482 10368
rect 18546 10304 18562 10368
rect 18626 10304 18634 10368
rect 18314 9280 18634 10304
rect 18314 9216 18322 9280
rect 18386 9216 18402 9280
rect 18466 9216 18482 9280
rect 18546 9216 18562 9280
rect 18626 9216 18634 9280
rect 18314 8192 18634 9216
rect 18314 8128 18322 8192
rect 18386 8128 18402 8192
rect 18466 8128 18482 8192
rect 18546 8128 18562 8192
rect 18626 8128 18634 8192
rect 18314 7104 18634 8128
rect 18314 7040 18322 7104
rect 18386 7040 18402 7104
rect 18466 7040 18482 7104
rect 18546 7040 18562 7104
rect 18626 7040 18634 7104
rect 18314 6016 18634 7040
rect 18314 5952 18322 6016
rect 18386 5952 18402 6016
rect 18466 5952 18482 6016
rect 18546 5952 18562 6016
rect 18626 5952 18634 6016
rect 18314 4928 18634 5952
rect 18314 4864 18322 4928
rect 18386 4864 18402 4928
rect 18466 4864 18482 4928
rect 18546 4864 18562 4928
rect 18626 4864 18634 4928
rect 18314 3840 18634 4864
rect 18314 3776 18322 3840
rect 18386 3776 18402 3840
rect 18466 3776 18482 3840
rect 18546 3776 18562 3840
rect 18626 3776 18634 3840
rect 18314 2752 18634 3776
rect 18314 2688 18322 2752
rect 18386 2688 18402 2752
rect 18466 2688 18482 2752
rect 18546 2688 18562 2752
rect 18626 2688 18634 2752
rect 18314 2128 18634 2688
rect 21788 27232 22108 27792
rect 21788 27168 21796 27232
rect 21860 27168 21876 27232
rect 21940 27168 21956 27232
rect 22020 27168 22036 27232
rect 22100 27168 22108 27232
rect 21788 26144 22108 27168
rect 21788 26080 21796 26144
rect 21860 26080 21876 26144
rect 21940 26080 21956 26144
rect 22020 26080 22036 26144
rect 22100 26080 22108 26144
rect 21788 25056 22108 26080
rect 21788 24992 21796 25056
rect 21860 24992 21876 25056
rect 21940 24992 21956 25056
rect 22020 24992 22036 25056
rect 22100 24992 22108 25056
rect 21788 23968 22108 24992
rect 21788 23904 21796 23968
rect 21860 23904 21876 23968
rect 21940 23904 21956 23968
rect 22020 23904 22036 23968
rect 22100 23904 22108 23968
rect 21788 22880 22108 23904
rect 21788 22816 21796 22880
rect 21860 22816 21876 22880
rect 21940 22816 21956 22880
rect 22020 22816 22036 22880
rect 22100 22816 22108 22880
rect 21788 21792 22108 22816
rect 21788 21728 21796 21792
rect 21860 21728 21876 21792
rect 21940 21728 21956 21792
rect 22020 21728 22036 21792
rect 22100 21728 22108 21792
rect 21788 20704 22108 21728
rect 21788 20640 21796 20704
rect 21860 20640 21876 20704
rect 21940 20640 21956 20704
rect 22020 20640 22036 20704
rect 22100 20640 22108 20704
rect 21788 19616 22108 20640
rect 21788 19552 21796 19616
rect 21860 19552 21876 19616
rect 21940 19552 21956 19616
rect 22020 19552 22036 19616
rect 22100 19552 22108 19616
rect 21788 18528 22108 19552
rect 21788 18464 21796 18528
rect 21860 18464 21876 18528
rect 21940 18464 21956 18528
rect 22020 18464 22036 18528
rect 22100 18464 22108 18528
rect 21788 17440 22108 18464
rect 21788 17376 21796 17440
rect 21860 17376 21876 17440
rect 21940 17376 21956 17440
rect 22020 17376 22036 17440
rect 22100 17376 22108 17440
rect 21788 16352 22108 17376
rect 21788 16288 21796 16352
rect 21860 16288 21876 16352
rect 21940 16288 21956 16352
rect 22020 16288 22036 16352
rect 22100 16288 22108 16352
rect 21788 15264 22108 16288
rect 21788 15200 21796 15264
rect 21860 15200 21876 15264
rect 21940 15200 21956 15264
rect 22020 15200 22036 15264
rect 22100 15200 22108 15264
rect 21788 14176 22108 15200
rect 21788 14112 21796 14176
rect 21860 14112 21876 14176
rect 21940 14112 21956 14176
rect 22020 14112 22036 14176
rect 22100 14112 22108 14176
rect 21788 13088 22108 14112
rect 21788 13024 21796 13088
rect 21860 13024 21876 13088
rect 21940 13024 21956 13088
rect 22020 13024 22036 13088
rect 22100 13024 22108 13088
rect 21788 12000 22108 13024
rect 21788 11936 21796 12000
rect 21860 11936 21876 12000
rect 21940 11936 21956 12000
rect 22020 11936 22036 12000
rect 22100 11936 22108 12000
rect 21788 10912 22108 11936
rect 21788 10848 21796 10912
rect 21860 10848 21876 10912
rect 21940 10848 21956 10912
rect 22020 10848 22036 10912
rect 22100 10848 22108 10912
rect 21788 9824 22108 10848
rect 21788 9760 21796 9824
rect 21860 9760 21876 9824
rect 21940 9760 21956 9824
rect 22020 9760 22036 9824
rect 22100 9760 22108 9824
rect 21788 8736 22108 9760
rect 21788 8672 21796 8736
rect 21860 8672 21876 8736
rect 21940 8672 21956 8736
rect 22020 8672 22036 8736
rect 22100 8672 22108 8736
rect 21788 7648 22108 8672
rect 21788 7584 21796 7648
rect 21860 7584 21876 7648
rect 21940 7584 21956 7648
rect 22020 7584 22036 7648
rect 22100 7584 22108 7648
rect 21788 6560 22108 7584
rect 21788 6496 21796 6560
rect 21860 6496 21876 6560
rect 21940 6496 21956 6560
rect 22020 6496 22036 6560
rect 22100 6496 22108 6560
rect 21788 5472 22108 6496
rect 21788 5408 21796 5472
rect 21860 5408 21876 5472
rect 21940 5408 21956 5472
rect 22020 5408 22036 5472
rect 22100 5408 22108 5472
rect 21788 4384 22108 5408
rect 21788 4320 21796 4384
rect 21860 4320 21876 4384
rect 21940 4320 21956 4384
rect 22020 4320 22036 4384
rect 22100 4320 22108 4384
rect 21788 3296 22108 4320
rect 21788 3232 21796 3296
rect 21860 3232 21876 3296
rect 21940 3232 21956 3296
rect 22020 3232 22036 3296
rect 22100 3232 22108 3296
rect 21788 2208 22108 3232
rect 21788 2144 21796 2208
rect 21860 2144 21876 2208
rect 21940 2144 21956 2208
rect 22020 2144 22036 2208
rect 22100 2144 22108 2208
rect 21788 2128 22108 2144
rect 25262 27776 25582 27792
rect 25262 27712 25270 27776
rect 25334 27712 25350 27776
rect 25414 27712 25430 27776
rect 25494 27712 25510 27776
rect 25574 27712 25582 27776
rect 25262 26688 25582 27712
rect 25262 26624 25270 26688
rect 25334 26624 25350 26688
rect 25414 26624 25430 26688
rect 25494 26624 25510 26688
rect 25574 26624 25582 26688
rect 25262 25600 25582 26624
rect 25262 25536 25270 25600
rect 25334 25536 25350 25600
rect 25414 25536 25430 25600
rect 25494 25536 25510 25600
rect 25574 25536 25582 25600
rect 25262 24512 25582 25536
rect 25262 24448 25270 24512
rect 25334 24448 25350 24512
rect 25414 24448 25430 24512
rect 25494 24448 25510 24512
rect 25574 24448 25582 24512
rect 25262 23424 25582 24448
rect 25262 23360 25270 23424
rect 25334 23360 25350 23424
rect 25414 23360 25430 23424
rect 25494 23360 25510 23424
rect 25574 23360 25582 23424
rect 25262 22336 25582 23360
rect 25262 22272 25270 22336
rect 25334 22272 25350 22336
rect 25414 22272 25430 22336
rect 25494 22272 25510 22336
rect 25574 22272 25582 22336
rect 25262 21248 25582 22272
rect 25262 21184 25270 21248
rect 25334 21184 25350 21248
rect 25414 21184 25430 21248
rect 25494 21184 25510 21248
rect 25574 21184 25582 21248
rect 25262 20160 25582 21184
rect 25262 20096 25270 20160
rect 25334 20096 25350 20160
rect 25414 20096 25430 20160
rect 25494 20096 25510 20160
rect 25574 20096 25582 20160
rect 25262 19072 25582 20096
rect 25262 19008 25270 19072
rect 25334 19008 25350 19072
rect 25414 19008 25430 19072
rect 25494 19008 25510 19072
rect 25574 19008 25582 19072
rect 25262 17984 25582 19008
rect 25262 17920 25270 17984
rect 25334 17920 25350 17984
rect 25414 17920 25430 17984
rect 25494 17920 25510 17984
rect 25574 17920 25582 17984
rect 25262 16896 25582 17920
rect 25262 16832 25270 16896
rect 25334 16832 25350 16896
rect 25414 16832 25430 16896
rect 25494 16832 25510 16896
rect 25574 16832 25582 16896
rect 25262 15808 25582 16832
rect 25262 15744 25270 15808
rect 25334 15744 25350 15808
rect 25414 15744 25430 15808
rect 25494 15744 25510 15808
rect 25574 15744 25582 15808
rect 25262 14720 25582 15744
rect 25262 14656 25270 14720
rect 25334 14656 25350 14720
rect 25414 14656 25430 14720
rect 25494 14656 25510 14720
rect 25574 14656 25582 14720
rect 25262 13632 25582 14656
rect 25262 13568 25270 13632
rect 25334 13568 25350 13632
rect 25414 13568 25430 13632
rect 25494 13568 25510 13632
rect 25574 13568 25582 13632
rect 25262 12544 25582 13568
rect 25262 12480 25270 12544
rect 25334 12480 25350 12544
rect 25414 12480 25430 12544
rect 25494 12480 25510 12544
rect 25574 12480 25582 12544
rect 25262 11456 25582 12480
rect 25262 11392 25270 11456
rect 25334 11392 25350 11456
rect 25414 11392 25430 11456
rect 25494 11392 25510 11456
rect 25574 11392 25582 11456
rect 25262 10368 25582 11392
rect 25262 10304 25270 10368
rect 25334 10304 25350 10368
rect 25414 10304 25430 10368
rect 25494 10304 25510 10368
rect 25574 10304 25582 10368
rect 25262 9280 25582 10304
rect 25262 9216 25270 9280
rect 25334 9216 25350 9280
rect 25414 9216 25430 9280
rect 25494 9216 25510 9280
rect 25574 9216 25582 9280
rect 25262 8192 25582 9216
rect 25262 8128 25270 8192
rect 25334 8128 25350 8192
rect 25414 8128 25430 8192
rect 25494 8128 25510 8192
rect 25574 8128 25582 8192
rect 25262 7104 25582 8128
rect 25262 7040 25270 7104
rect 25334 7040 25350 7104
rect 25414 7040 25430 7104
rect 25494 7040 25510 7104
rect 25574 7040 25582 7104
rect 25262 6016 25582 7040
rect 25262 5952 25270 6016
rect 25334 5952 25350 6016
rect 25414 5952 25430 6016
rect 25494 5952 25510 6016
rect 25574 5952 25582 6016
rect 25262 4928 25582 5952
rect 25262 4864 25270 4928
rect 25334 4864 25350 4928
rect 25414 4864 25430 4928
rect 25494 4864 25510 4928
rect 25574 4864 25582 4928
rect 25262 3840 25582 4864
rect 25262 3776 25270 3840
rect 25334 3776 25350 3840
rect 25414 3776 25430 3840
rect 25494 3776 25510 3840
rect 25574 3776 25582 3840
rect 25262 2752 25582 3776
rect 25262 2688 25270 2752
rect 25334 2688 25350 2752
rect 25414 2688 25430 2752
rect 25494 2688 25510 2752
rect 25574 2688 25582 2752
rect 25262 2128 25582 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A0 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7636 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A0
timestamp 1649977179
transform 1 0 15272 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__A
timestamp 1649977179
transform -1 0 17112 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A
timestamp 1649977179
transform 1 0 5244 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__A
timestamp 1649977179
transform -1 0 1932 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A
timestamp 1649977179
transform 1 0 3956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1649977179
transform 1 0 17204 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1649977179
transform -1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A
timestamp 1649977179
transform -1 0 3772 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1649977179
transform -1 0 6256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 27600 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 17756 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 22908 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_233 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22540 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1649977179
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1649977179
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1649977179
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_293
timestamp 1649977179
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_36
timestamp 1649977179
transform 1 0 4416 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1649977179
transform 1 0 5244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_62
timestamp 1649977179
transform 1 0 6808 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_74
timestamp 1649977179
transform 1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_97
timestamp 1649977179
transform 1 0 10028 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_143
timestamp 1649977179
transform 1 0 14260 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_147
timestamp 1649977179
transform 1 0 14628 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_154
timestamp 1649977179
transform 1 0 15272 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1649977179
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1649977179
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1649977179
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1649977179
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1649977179
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1649977179
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_293
timestamp 1649977179
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_10
timestamp 1649977179
transform 1 0 2024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_17
timestamp 1649977179
transform 1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1649977179
transform 1 0 5796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75
timestamp 1649977179
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_88
timestamp 1649977179
transform 1 0 9200 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_100
timestamp 1649977179
transform 1 0 10304 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_161
timestamp 1649977179
transform 1 0 15916 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1649977179
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_289
timestamp 1649977179
transform 1 0 27692 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_297
timestamp 1649977179
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1649977179
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_30
timestamp 1649977179
transform 1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_42
timestamp 1649977179
transform 1 0 4968 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1649977179
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_77
timestamp 1649977179
transform 1 0 8188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_89
timestamp 1649977179
transform 1 0 9292 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_101
timestamp 1649977179
transform 1 0 10396 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1649977179
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_133
timestamp 1649977179
transform 1 0 13340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_145
timestamp 1649977179
transform 1 0 14444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_157
timestamp 1649977179
transform 1 0 15548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp 1649977179
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1649977179
transform 1 0 4048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1649977179
transform 1 0 4416 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_40
timestamp 1649977179
transform 1 0 4784 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_52
timestamp 1649977179
transform 1 0 5888 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_56
timestamp 1649977179
transform 1 0 6256 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_120
timestamp 1649977179
transform 1 0 12144 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_132
timestamp 1649977179
transform 1 0 13248 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_144
timestamp 1649977179
transform 1 0 14352 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_151
timestamp 1649977179
transform 1 0 14996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_163
timestamp 1649977179
transform 1 0 16100 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_168
timestamp 1649977179
transform 1 0 16560 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_174
timestamp 1649977179
transform 1 0 17112 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_186
timestamp 1649977179
transform 1 0 18216 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1649977179
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_206
timestamp 1649977179
transform 1 0 20056 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_218
timestamp 1649977179
transform 1 0 21160 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_230
timestamp 1649977179
transform 1 0 22264 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_242
timestamp 1649977179
transform 1 0 23368 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1649977179
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1649977179
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_14
timestamp 1649977179
transform 1 0 2392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1649977179
transform 1 0 4600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_48
timestamp 1649977179
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_64
timestamp 1649977179
transform 1 0 6992 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_72
timestamp 1649977179
transform 1 0 7728 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_100
timestamp 1649977179
transform 1 0 10304 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_116
timestamp 1649977179
transform 1 0 11776 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_128
timestamp 1649977179
transform 1 0 12880 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_139
timestamp 1649977179
transform 1 0 13892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_151
timestamp 1649977179
transform 1 0 14996 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_163
timestamp 1649977179
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_63
timestamp 1649977179
transform 1 0 6900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1649977179
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1649977179
transform 1 0 9200 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_92
timestamp 1649977179
transform 1 0 9568 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_113
timestamp 1649977179
transform 1 0 11500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_125
timestamp 1649977179
transform 1 0 12604 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1649977179
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_145
timestamp 1649977179
transform 1 0 14444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_164
timestamp 1649977179
transform 1 0 16192 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_176
timestamp 1649977179
transform 1 0 17296 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_188
timestamp 1649977179
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_297
timestamp 1649977179
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1649977179
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_30
timestamp 1649977179
transform 1 0 3864 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_41
timestamp 1649977179
transform 1 0 4876 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1649977179
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_77
timestamp 1649977179
transform 1 0 8188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_101
timestamp 1649977179
transform 1 0 10396 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1649977179
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_116
timestamp 1649977179
transform 1 0 11776 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_124
timestamp 1649977179
transform 1 0 12512 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_133
timestamp 1649977179
transform 1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_143
timestamp 1649977179
transform 1 0 14260 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_151
timestamp 1649977179
transform 1 0 14996 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_163
timestamp 1649977179
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_9
timestamp 1649977179
transform 1 0 1932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_16
timestamp 1649977179
transform 1 0 2576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1649977179
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_105
timestamp 1649977179
transform 1 0 10764 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_126
timestamp 1649977179
transform 1 0 12696 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1649977179
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_147
timestamp 1649977179
transform 1 0 14628 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_159
timestamp 1649977179
transform 1 0 15732 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_172
timestamp 1649977179
transform 1 0 16928 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_184
timestamp 1649977179
transform 1 0 18032 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_297
timestamp 1649977179
transform 1 0 28428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_12
timestamp 1649977179
transform 1 0 2208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_36
timestamp 1649977179
transform 1 0 4416 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_45
timestamp 1649977179
transform 1 0 5244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_87
timestamp 1649977179
transform 1 0 9108 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_136
timestamp 1649977179
transform 1 0 13616 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_143
timestamp 1649977179
transform 1 0 14260 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_150
timestamp 1649977179
transform 1 0 14904 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp 1649977179
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1649977179
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_32
timestamp 1649977179
transform 1 0 4048 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_44
timestamp 1649977179
transform 1 0 5152 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_52
timestamp 1649977179
transform 1 0 5888 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_56
timestamp 1649977179
transform 1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1649977179
transform 1 0 9660 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_123
timestamp 1649977179
transform 1 0 12420 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_131
timestamp 1649977179
transform 1 0 13156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_147
timestamp 1649977179
transform 1 0 14628 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_158
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_166
timestamp 1649977179
transform 1 0 16376 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_171
timestamp 1649977179
transform 1 0 16836 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_297
timestamp 1649977179
transform 1 0 28428 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_43
timestamp 1649977179
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_68
timestamp 1649977179
transform 1 0 7360 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_80
timestamp 1649977179
transform 1 0 8464 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1649977179
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_116
timestamp 1649977179
transform 1 0 11776 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_128
timestamp 1649977179
transform 1 0 12880 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_136
timestamp 1649977179
transform 1 0 13616 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_142
timestamp 1649977179
transform 1 0 14168 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_154
timestamp 1649977179
transform 1 0 15272 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_73
timestamp 1649977179
transform 1 0 7820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1649977179
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_100
timestamp 1649977179
transform 1 0 10304 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_112
timestamp 1649977179
transform 1 0 11408 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_124
timestamp 1649977179
transform 1 0 12512 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_146
timestamp 1649977179
transform 1 0 14536 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_158
timestamp 1649977179
transform 1 0 15640 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_170
timestamp 1649977179
transform 1 0 16744 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_182
timestamp 1649977179
transform 1 0 17848 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1649977179
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_297
timestamp 1649977179
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_80
timestamp 1649977179
transform 1 0 8464 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_92
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_104
timestamp 1649977179
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_133
timestamp 1649977179
transform 1 0 13340 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_139
timestamp 1649977179
transform 1 0 13892 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_145
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_171
timestamp 1649977179
transform 1 0 16836 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_183
timestamp 1649977179
transform 1 0 17940 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_191
timestamp 1649977179
transform 1 0 18676 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_196
timestamp 1649977179
transform 1 0 19136 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_203
timestamp 1649977179
transform 1 0 19780 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1649977179
transform 1 0 20884 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_76
timestamp 1649977179
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_120
timestamp 1649977179
transform 1 0 12144 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_132
timestamp 1649977179
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_148
timestamp 1649977179
transform 1 0 14720 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_160
timestamp 1649977179
transform 1 0 15824 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_172
timestamp 1649977179
transform 1 0 16928 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_184
timestamp 1649977179
transform 1 0 18032 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp 1649977179
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1649977179
transform 1 0 1748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_28
timestamp 1649977179
transform 1 0 3680 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_78
timestamp 1649977179
transform 1 0 8280 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_84
timestamp 1649977179
transform 1 0 8832 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_106
timestamp 1649977179
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_133
timestamp 1649977179
transform 1 0 13340 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_145
timestamp 1649977179
transform 1 0 14444 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_152
timestamp 1649977179
transform 1 0 15088 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1649977179
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1649977179
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_51
timestamp 1649977179
transform 1 0 5796 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_63
timestamp 1649977179
transform 1 0 6900 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_75
timestamp 1649977179
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_101
timestamp 1649977179
transform 1 0 10396 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_122
timestamp 1649977179
transform 1 0 12328 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_134
timestamp 1649977179
transform 1 0 13432 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_147
timestamp 1649977179
transform 1 0 14628 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_151
timestamp 1649977179
transform 1 0 14996 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_163
timestamp 1649977179
transform 1 0 16100 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_175
timestamp 1649977179
transform 1 0 17204 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_187
timestamp 1649977179
transform 1 0 18308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1649977179
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_35
timestamp 1649977179
transform 1 0 4324 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_41
timestamp 1649977179
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1649977179
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_101
timestamp 1649977179
transform 1 0 10396 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1649977179
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_116
timestamp 1649977179
transform 1 0 11776 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_128
timestamp 1649977179
transform 1 0 12880 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_140
timestamp 1649977179
transform 1 0 13984 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_152
timestamp 1649977179
transform 1 0 15088 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_45
timestamp 1649977179
transform 1 0 5244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_57
timestamp 1649977179
transform 1 0 6348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_69
timestamp 1649977179
transform 1 0 7452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp 1649977179
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_150
timestamp 1649977179
transform 1 0 14904 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_156
timestamp 1649977179
transform 1 0 15456 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_168
timestamp 1649977179
transform 1 0 16560 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_180
timestamp 1649977179
transform 1 0 17664 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp 1649977179
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_29
timestamp 1649977179
transform 1 0 3772 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_36
timestamp 1649977179
transform 1 0 4416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_43
timestamp 1649977179
transform 1 0 5060 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1649977179
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_61
timestamp 1649977179
transform 1 0 6716 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_65
timestamp 1649977179
transform 1 0 7084 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_72
timestamp 1649977179
transform 1 0 7728 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_84
timestamp 1649977179
transform 1 0 8832 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_119
timestamp 1649977179
transform 1 0 12052 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_131
timestamp 1649977179
transform 1 0 13156 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_142
timestamp 1649977179
transform 1 0 14168 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_150
timestamp 1649977179
transform 1 0 14904 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1649977179
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_9
timestamp 1649977179
transform 1 0 1932 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1649977179
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_37
timestamp 1649977179
transform 1 0 4508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_44
timestamp 1649977179
transform 1 0 5152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_51
timestamp 1649977179
transform 1 0 5796 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_64
timestamp 1649977179
transform 1 0 6992 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_75
timestamp 1649977179
transform 1 0 8004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_89
timestamp 1649977179
transform 1 0 9292 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_98
timestamp 1649977179
transform 1 0 10120 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_107
timestamp 1649977179
transform 1 0 10948 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_114
timestamp 1649977179
transform 1 0 11592 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_127
timestamp 1649977179
transform 1 0 12788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_146
timestamp 1649977179
transform 1 0 14536 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_154
timestamp 1649977179
transform 1 0 15272 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_166
timestamp 1649977179
transform 1 0 16376 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_178
timestamp 1649977179
transform 1 0 17480 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1649977179
transform 1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1649977179
transform 1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_12
timestamp 1649977179
transform 1 0 2208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_23
timestamp 1649977179
transform 1 0 3220 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_37
timestamp 1649977179
transform 1 0 4508 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1649977179
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_61
timestamp 1649977179
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_71
timestamp 1649977179
transform 1 0 7636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_78
timestamp 1649977179
transform 1 0 8280 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_82
timestamp 1649977179
transform 1 0 8648 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_90
timestamp 1649977179
transform 1 0 9384 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_94
timestamp 1649977179
transform 1 0 9752 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_102
timestamp 1649977179
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1649977179
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_135
timestamp 1649977179
transform 1 0 13524 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_142
timestamp 1649977179
transform 1 0 14168 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_154
timestamp 1649977179
transform 1 0 15272 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1649977179
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_17
timestamp 1649977179
transform 1 0 2668 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1649977179
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_33
timestamp 1649977179
transform 1 0 4140 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_45
timestamp 1649977179
transform 1 0 5244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_57
timestamp 1649977179
transform 1 0 6348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_61
timestamp 1649977179
transform 1 0 6716 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_73
timestamp 1649977179
transform 1 0 7820 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1649977179
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_106
timestamp 1649977179
transform 1 0 10856 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_117
timestamp 1649977179
transform 1 0 11868 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_124
timestamp 1649977179
transform 1 0 12512 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1649977179
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_297
timestamp 1649977179
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_14
timestamp 1649977179
transform 1 0 2392 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_26
timestamp 1649977179
transform 1 0 3496 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_34
timestamp 1649977179
transform 1 0 4232 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_42
timestamp 1649977179
transform 1 0 4968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_60
timestamp 1649977179
transform 1 0 6624 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_68
timestamp 1649977179
transform 1 0 7360 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_73
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_85
timestamp 1649977179
transform 1 0 8924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_97
timestamp 1649977179
transform 1 0 10028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_126
timestamp 1649977179
transform 1 0 12696 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_138
timestamp 1649977179
transform 1 0 13800 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_150
timestamp 1649977179
transform 1 0 14904 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_162
timestamp 1649977179
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_45
timestamp 1649977179
transform 1 0 5244 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_54
timestamp 1649977179
transform 1 0 6072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_61
timestamp 1649977179
transform 1 0 6716 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_70
timestamp 1649977179
transform 1 0 7544 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1649977179
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_92
timestamp 1649977179
transform 1 0 9568 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_104
timestamp 1649977179
transform 1 0 10672 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_112
timestamp 1649977179
transform 1 0 11408 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_120
timestamp 1649977179
transform 1 0 12144 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_126
timestamp 1649977179
transform 1 0 12696 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1649977179
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_31
timestamp 1649977179
transform 1 0 3956 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_46
timestamp 1649977179
transform 1 0 5336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1649977179
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_61
timestamp 1649977179
transform 1 0 6716 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_78
timestamp 1649977179
transform 1 0 8280 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_82
timestamp 1649977179
transform 1 0 8648 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_90
timestamp 1649977179
transform 1 0 9384 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_102
timestamp 1649977179
transform 1 0 10488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1649977179
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_121
timestamp 1649977179
transform 1 0 12236 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_133
timestamp 1649977179
transform 1 0 13340 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_145
timestamp 1649977179
transform 1 0 14444 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_157
timestamp 1649977179
transform 1 0 15548 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1649977179
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_37
timestamp 1649977179
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_49
timestamp 1649977179
transform 1 0 5612 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_61
timestamp 1649977179
transform 1 0 6716 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_66
timestamp 1649977179
transform 1 0 7176 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1649977179
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_94
timestamp 1649977179
transform 1 0 9752 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_103
timestamp 1649977179
transform 1 0 10580 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_117
timestamp 1649977179
transform 1 0 11868 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_129
timestamp 1649977179
transform 1 0 12972 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1649977179
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_297
timestamp 1649977179
transform 1 0 28428 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_35
timestamp 1649977179
transform 1 0 4324 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_44
timestamp 1649977179
transform 1 0 5152 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_76
timestamp 1649977179
transform 1 0 8096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_80
timestamp 1649977179
transform 1 0 8464 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_88
timestamp 1649977179
transform 1 0 9200 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_100
timestamp 1649977179
transform 1 0 10304 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_285
timestamp 1649977179
transform 1 0 27324 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_288
timestamp 1649977179
transform 1 0 27600 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_295
timestamp 1649977179
transform 1 0 28244 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_289
timestamp 1649977179
transform 1 0 27692 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_297
timestamp 1649977179
transform 1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_297
timestamp 1649977179
transform 1 0 28428 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1649977179
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_31
timestamp 1649977179
transform 1 0 3956 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_43
timestamp 1649977179
transform 1 0 5060 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_55
timestamp 1649977179
transform 1 0 6164 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_67
timestamp 1649977179
transform 1 0 7268 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp 1649977179
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp 1649977179
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_23
timestamp 1649977179
transform 1 0 3220 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_33
timestamp 1649977179
transform 1 0 4140 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_45
timestamp 1649977179
transform 1 0 5244 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1649977179
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp 1649977179
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1649977179
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_297
timestamp 1649977179
transform 1 0 28428 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1649977179
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1649977179
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1649977179
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_289
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_297
timestamp 1649977179
transform 1 0 28428 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1649977179
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1649977179
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1649977179
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1649977179
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1649977179
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1649977179
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1649977179
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1649977179
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1649977179
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1649977179
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1649977179
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_289
timestamp 1649977179
transform 1 0 27692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_297
timestamp 1649977179
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_7
timestamp 1649977179
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_19
timestamp 1649977179
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_31
timestamp 1649977179
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_43
timestamp 1649977179
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1649977179
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1649977179
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1649977179
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1649977179
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1649977179
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1649977179
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_289
timestamp 1649977179
transform 1 0 27692 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp 1649977179
transform 1 0 28428 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1649977179
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1649977179
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1649977179
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1649977179
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1649977179
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1649977179
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1649977179
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1649977179
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_289
timestamp 1649977179
transform 1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_297
timestamp 1649977179
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1649977179
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1649977179
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1649977179
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1649977179
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1649977179
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1649977179
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1649977179
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1649977179
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_57
timestamp 1649977179
transform 1 0 6348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_69
timestamp 1649977179
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1649977179
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_113
timestamp 1649977179
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_125
timestamp 1649977179
transform 1 0 12604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1649977179
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_169
timestamp 1649977179
transform 1 0 16652 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_177
timestamp 1649977179
transform 1 0 17388 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_181
timestamp 1649977179
transform 1 0 17756 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_188
timestamp 1649977179
transform 1 0 18400 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_221
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_225
timestamp 1649977179
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_237
timestamp 1649977179
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1649977179
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1649977179
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_277
timestamp 1649977179
transform 1 0 26588 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_281
timestamp 1649977179
transform 1 0 26956 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_293
timestamp 1649977179
transform 1 0 28060 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _142_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _143_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13984 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _144_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _145_
timestamp 1649977179
transform 1 0 12788 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _146_
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _147_
timestamp 1649977179
transform 1 0 14628 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _148_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _149_
timestamp 1649977179
transform 1 0 6348 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _150_
timestamp 1649977179
transform 1 0 4968 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _151_
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _152_
timestamp 1649977179
transform -1 0 14536 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _153_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12604 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _154_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _155_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6164 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _156_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4968 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _157_
timestamp 1649977179
transform -1 0 7636 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1649977179
transform -1 0 7728 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _159_
timestamp 1649977179
transform 1 0 11960 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1649977179
transform 1 0 11776 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _161_
timestamp 1649977179
transform -1 0 14904 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12512 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _164_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7820 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _165_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9844 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _166_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9200 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _167_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9660 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _168_
timestamp 1649977179
transform -1 0 13524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _169_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11868 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _170_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11316 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1649977179
transform -1 0 7544 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _172_
timestamp 1649977179
transform 1 0 8740 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1649977179
transform 1 0 8004 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1649977179
transform -1 0 7176 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1649977179
transform -1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1649977179
transform -1 0 6716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _177_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6072 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _178_
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _179_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10580 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _180_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9108 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _181_
timestamp 1649977179
transform -1 0 8096 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _182_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8372 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _183_
timestamp 1649977179
transform -1 0 10948 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _184_
timestamp 1649977179
transform 1 0 8740 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _185_
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _186_
timestamp 1649977179
transform 1 0 6440 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _187_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11684 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _188_
timestamp 1649977179
transform 1 0 12052 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _189_
timestamp 1649977179
transform 1 0 12788 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1649977179
transform 1 0 11316 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _191_
timestamp 1649977179
transform 1 0 5244 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _192_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14168 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _193_
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _194_
timestamp 1649977179
transform -1 0 3956 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _195_
timestamp 1649977179
transform 1 0 2576 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _196_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _197_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4140 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _198_
timestamp 1649977179
transform 1 0 2116 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _199_
timestamp 1649977179
transform -1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _200_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _201_
timestamp 1649977179
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _202_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1656 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _203_
timestamp 1649977179
transform 1 0 3036 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _204_
timestamp 1649977179
transform -1 0 4968 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _205_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _206_
timestamp 1649977179
transform 1 0 4600 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _207_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4784 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _208_
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _209_
timestamp 1649977179
transform 1 0 14996 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _210_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15272 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1649977179
transform -1 0 8464 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _212_
timestamp 1649977179
transform -1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _213_
timestamp 1649977179
transform -1 0 7084 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1649977179
transform -1 0 8004 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1649977179
transform 1 0 9384 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _216_
timestamp 1649977179
transform 1 0 14628 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1649977179
transform -1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1649977179
transform -1 0 19136 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1649977179
transform -1 0 13616 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1649977179
transform -1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1649977179
transform 1 0 19504 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _222_
timestamp 1649977179
transform -1 0 15180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1649977179
transform -1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 1649977179
transform -1 0 14628 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1649977179
transform -1 0 4784 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1649977179
transform -1 0 15272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1649977179
transform 1 0 15916 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _228_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16376 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1649977179
transform 1 0 2760 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1649977179
transform -1 0 16560 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1649977179
transform -1 0 4876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1649977179
transform -1 0 3220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1649977179
transform -1 0 3588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _234_
timestamp 1649977179
transform -1 0 14444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1649977179
transform -1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1649977179
transform 1 0 19780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1649977179
transform -1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1649977179
transform -1 0 13616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1649977179
transform -1 0 14996 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _240_
timestamp 1649977179
transform -1 0 16836 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1649977179
transform -1 0 14904 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1649977179
transform -1 0 14168 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1649977179
transform -1 0 13616 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1649977179
transform -1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1649977179
transform -1 0 14260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _246_
timestamp 1649977179
transform -1 0 12144 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1649977179
transform -1 0 5796 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1649977179
transform 1 0 9016 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1649977179
transform -1 0 14168 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1649977179
transform 1 0 14720 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1649977179
transform -1 0 14720 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _252_
timestamp 1649977179
transform 1 0 4140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1649977179
transform -1 0 5060 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1649977179
transform 1 0 5428 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1649977179
transform -1 0 5152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1649977179
transform -1 0 5244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1649977179
transform -1 0 4416 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_2  _258_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _259_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10856 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _260_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6164 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _261_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _262_
timestamp 1649977179
transform 1 0 10488 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _263__31 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _263_
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _264__30
timestamp 1649977179
transform -1 0 7360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _264_
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _265__29
timestamp 1649977179
transform -1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _265_
timestamp 1649977179
transform 1 0 4140 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _266__28
timestamp 1649977179
transform -1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _266_
timestamp 1649977179
transform 1 0 8188 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _267__27
timestamp 1649977179
transform -1 0 6992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _267_
timestamp 1649977179
transform 1 0 6348 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _268_
timestamp 1649977179
transform 1 0 3956 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _268__26
timestamp 1649977179
transform -1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _269_
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _269__25
timestamp 1649977179
transform -1 0 11040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _270_
timestamp 1649977179
transform 1 0 2024 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _270__24
timestamp 1649977179
transform -1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _271_
timestamp 1649977179
transform 1 0 6164 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _271__23
timestamp 1649977179
transform -1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _272__22
timestamp 1649977179
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _272_
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _273__21
timestamp 1649977179
transform -1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _273_
timestamp 1649977179
transform 1 0 2024 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _274__20
timestamp 1649977179
transform -1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _274_
timestamp 1649977179
transform 1 0 1472 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _275_
timestamp 1649977179
transform 1 0 3220 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _275__19
timestamp 1649977179
transform -1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _276__18
timestamp 1649977179
transform -1 0 2392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _276_
timestamp 1649977179
transform 1 0 1472 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _277_
timestamp 1649977179
transform 1 0 1472 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _277__17
timestamp 1649977179
transform -1 0 2208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _278__16
timestamp 1649977179
transform -1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _278_
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _279_
timestamp 1649977179
transform 1 0 2760 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _279__15
timestamp 1649977179
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _280_
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _280__14
timestamp 1649977179
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _281_
timestamp 1649977179
transform 1 0 9660 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _281__13
timestamp 1649977179
transform -1 0 10304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _282_
timestamp 1649977179
transform 1 0 10304 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _282__12
timestamp 1649977179
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _283_
timestamp 1649977179
transform 1 0 10856 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _283__11
timestamp 1649977179
transform -1 0 11776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _284__10
timestamp 1649977179
transform -1 0 10304 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _284_
timestamp 1649977179
transform 1 0 9200 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _285_
timestamp 1649977179
transform 1 0 9200 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _285__9
timestamp 1649977179
transform -1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _286__8
timestamp 1649977179
transform -1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _286_
timestamp 1649977179
transform 1 0 10304 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _287__7
timestamp 1649977179
transform -1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _287_
timestamp 1649977179
transform 1 0 10580 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _288__6
timestamp 1649977179
transform -1 0 4876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _288_
timestamp 1649977179
transform 1 0 4048 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _289__5
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _289_
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _290_
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _291_
timestamp 1649977179
transform 1 0 7820 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _292_
timestamp 1649977179
transform -1 0 8464 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _293_
timestamp 1649977179
transform 1 0 1472 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _294_
timestamp 1649977179
transform 1 0 1840 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _295_
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _296_
timestamp 1649977179
transform 1 0 1472 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _297_
timestamp 1649977179
transform 1 0 3956 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6716 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1649977179
transform -1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1649977179
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1649977179
transform 1 0 7820 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1649977179
transform 1 0 6624 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform 1 0 27968 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform 1 0 18124 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1649977179
transform -1 0 23644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1649977179
transform -1 0 1748 0 -1 25024
box -38 -48 406 592
<< labels >>
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 PWM_OUT
port 0 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 clk
port 1 nsew signal input
flabel metal3 s 29200 17008 30000 17128 0 FreeSans 480 0 0 0 decrease_duty
port 2 nsew signal input
flabel metal2 s 18050 29200 18106 30000 0 FreeSans 224 90 0 0 increase_duty
port 3 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 reset
port 4 nsew signal input
flabel metal4 s 4418 2128 4738 27792 0 FreeSans 1920 90 0 0 vccd1
port 5 nsew power bidirectional
flabel metal4 s 11366 2128 11686 27792 0 FreeSans 1920 90 0 0 vccd1
port 5 nsew power bidirectional
flabel metal4 s 18314 2128 18634 27792 0 FreeSans 1920 90 0 0 vccd1
port 5 nsew power bidirectional
flabel metal4 s 25262 2128 25582 27792 0 FreeSans 1920 90 0 0 vccd1
port 5 nsew power bidirectional
flabel metal4 s 7892 2128 8212 27792 0 FreeSans 1920 90 0 0 vssd1
port 6 nsew ground bidirectional
flabel metal4 s 14840 2128 15160 27792 0 FreeSans 1920 90 0 0 vssd1
port 6 nsew ground bidirectional
flabel metal4 s 21788 2128 22108 27792 0 FreeSans 1920 90 0 0 vssd1
port 6 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
